magic
tech sky130A
magscale 1 2
timestamp 1725111887
<< nwell >>
rect -1040 5660 16500 8780
rect 9590 160 16500 5660
<< pwell >>
rect 890 -560 8580 5060
rect 7580 -1870 16510 -1690
rect -1340 -4970 16510 -1870
<< mvpsubdiff >>
rect 960 4990 8510 5000
rect 960 4940 1120 4990
rect 8350 4940 8510 4990
rect 960 4930 8510 4940
rect 960 4880 1030 4930
rect 960 -370 970 4880
rect 1020 -370 1030 4880
rect 960 -410 1030 -370
rect 8440 4880 8510 4930
rect 8440 -370 8450 4880
rect 8500 -370 8510 4880
rect 8440 -410 8510 -370
rect 960 -420 8510 -410
rect 960 -470 1120 -420
rect 8350 -470 8510 -420
rect 960 -480 8510 -470
rect 7650 -1770 16440 -1760
rect 7650 -1820 7760 -1770
rect 16330 -1820 16440 -1770
rect 7650 -1830 16440 -1820
rect 7650 -1870 7720 -1830
rect -1270 -1950 7520 -1940
rect -1270 -2000 -1160 -1950
rect 7410 -2000 7520 -1950
rect -1270 -2010 7520 -2000
rect -1270 -2050 -1200 -2010
rect -1270 -4790 -1260 -2050
rect -1210 -4790 -1200 -2050
rect -1270 -4830 -1200 -4790
rect 7450 -2050 7520 -2010
rect 7450 -4790 7460 -2050
rect 7510 -4790 7520 -2050
rect 7450 -4830 7520 -4790
rect -1270 -4840 7520 -4830
rect -1270 -4890 -1160 -4840
rect 7410 -4890 7520 -4840
rect -1270 -4900 7520 -4890
rect 7650 -4790 7660 -1870
rect 7710 -4790 7720 -1870
rect 7650 -4830 7720 -4790
rect 16370 -1870 16440 -1830
rect 16370 -4790 16380 -1870
rect 16430 -4790 16440 -1870
rect 16370 -4830 16440 -4790
rect 7650 -4840 16440 -4830
rect 7650 -4890 7760 -4840
rect 16330 -4890 16440 -4840
rect 7650 -4900 16440 -4890
<< mvnsubdiff >>
rect -970 8700 16430 8710
rect -970 8650 -860 8700
rect 7650 8650 7810 8700
rect 16320 8650 16430 8700
rect -970 8640 16430 8650
rect -970 8600 -900 8640
rect -970 5880 -960 8600
rect -910 5880 -900 8600
rect -970 5840 -900 5880
rect 7690 8600 7770 8640
rect 7690 5880 7700 8600
rect 7760 5880 7770 8600
rect 7690 5840 7770 5880
rect 16360 8600 16430 8640
rect 16360 5880 16370 8600
rect 16420 5880 16430 8600
rect 16360 5840 16430 5880
rect -970 5830 16430 5840
rect -970 5780 -860 5830
rect 7650 5780 7810 5830
rect 16320 5780 16430 5830
rect -970 5770 16430 5780
rect 9660 5370 16080 5380
rect 9660 5320 9770 5370
rect 15970 5320 16080 5370
rect 9660 5310 16080 5320
rect 9660 5270 9730 5310
rect 9660 340 9670 5270
rect 9720 340 9730 5270
rect 9660 300 9730 340
rect 16010 5270 16080 5310
rect 16010 340 16020 5270
rect 16070 340 16080 5270
rect 16010 300 16080 340
rect 9660 290 16080 300
rect 9660 240 9770 290
rect 15970 240 16080 290
rect 9660 230 16080 240
<< mvpsubdiffcont >>
rect 1120 4940 8350 4990
rect 970 -370 1020 4880
rect 8450 -370 8500 4880
rect 1120 -470 8350 -420
rect 7760 -1820 16330 -1770
rect -1160 -2000 7410 -1950
rect -1260 -4790 -1210 -2050
rect 7460 -4790 7510 -2050
rect -1160 -4890 7410 -4840
rect 7660 -4790 7710 -1870
rect 16380 -4790 16430 -1870
rect 7760 -4890 16330 -4840
<< mvnsubdiffcont >>
rect -860 8650 7650 8700
rect 7810 8650 16320 8700
rect -960 5880 -910 8600
rect 7700 5880 7760 8600
rect 16370 5880 16420 8600
rect -860 5780 7650 5830
rect 7810 5780 16320 5830
rect 9770 5320 15970 5370
rect 9670 340 9720 5270
rect 16020 340 16070 5270
rect 9770 240 15970 290
<< locali >>
rect -960 8650 -860 8700
rect 7650 8650 7810 8700
rect 16320 8650 16420 8700
rect -960 8600 -910 8650
rect -960 5830 -910 5880
rect 7700 8600 7760 8650
rect 7700 5830 7760 5880
rect 16370 8600 16420 8650
rect 16370 5830 16420 5880
rect -960 5780 -860 5830
rect 7650 5780 7810 5830
rect 16320 5780 16420 5830
rect 9670 5320 9770 5370
rect 15970 5320 16070 5370
rect 9670 5270 9720 5320
rect 970 4940 1120 4990
rect 8350 4940 8500 4990
rect 970 4880 1020 4940
rect 970 -420 1020 -370
rect 8450 4880 8500 4940
rect 9670 290 9720 340
rect 16020 5270 16070 5320
rect 16020 290 16070 340
rect 9670 240 9770 290
rect 15970 240 16070 290
rect 8450 -420 8500 -370
rect 970 -470 1120 -420
rect 8350 -470 8500 -420
rect 7660 -1820 7760 -1770
rect 16330 -1820 16430 -1770
rect 7660 -1870 7710 -1820
rect -1260 -2000 -1160 -1950
rect 7410 -2000 7510 -1950
rect -1260 -2050 -1210 -2000
rect -1260 -4840 -1210 -4790
rect 7460 -2050 7510 -2000
rect 7460 -4840 7510 -4790
rect -1260 -4890 -1160 -4840
rect 7410 -4890 7510 -4840
rect 7660 -4840 7710 -4790
rect 16380 -1870 16430 -1820
rect 16380 -4840 16430 -4790
rect 7660 -4890 7760 -4840
rect 16330 -4890 16430 -4840
<< viali >>
rect -850 8650 7650 8700
rect 7810 8650 16320 8700
rect -960 5880 -910 8600
rect 7700 5880 7760 8600
rect 16370 5880 16420 8600
rect -860 5780 7650 5830
rect 7810 5780 16320 5830
rect 9770 5320 15970 5370
rect 1120 4940 8350 4990
rect 970 -370 1020 4880
rect 8450 -370 8500 4880
rect 9670 340 9720 5270
rect 16020 340 16070 5270
rect 9770 240 15970 290
rect 1120 -470 8350 -420
rect 14416 -1498 14450 -1148
rect 15874 -1498 15908 -1148
rect 14512 -1594 15812 -1560
rect 7760 -1820 16330 -1770
rect -1160 -2000 7410 -1950
rect -1260 -4790 -1210 -2050
rect 7460 -4790 7510 -2050
rect -1160 -4890 7410 -4840
rect 7660 -4790 7710 -1870
rect 16380 -4790 16430 -1870
rect 7760 -4890 16330 -4840
<< metal1 >>
rect -1490 8700 16500 9150
rect -1490 8650 -850 8700
rect 7650 8650 7810 8700
rect 16320 8650 16500 8700
rect -1490 8640 16500 8650
rect -1490 8600 -900 8640
rect -1490 5880 -960 8600
rect -910 5880 -900 8600
rect -1490 5840 -900 5880
rect 1585 8445 1662 8640
rect 1585 8343 1650 8445
rect 1585 6317 1662 8343
rect 1585 6215 1650 6317
rect 1585 5840 1662 6215
rect 1775 5840 1973 8640
rect 2086 8445 2163 8640
rect 2099 8343 2163 8445
rect 2086 6317 2163 8343
rect 2098 6215 2163 6317
rect 2086 5840 2163 6215
rect 2195 8445 2272 8640
rect 2385 8580 2583 8600
rect 2385 8460 2390 8580
rect 2570 8460 2583 8580
rect 2195 8343 2260 8445
rect 2195 6317 2272 8343
rect 2195 6215 2260 6317
rect 2195 6060 2272 6215
rect 2385 6200 2583 8460
rect 2696 8445 2773 8600
rect 2709 8343 2773 8445
rect 2696 6317 2773 8343
rect 2708 6215 2773 6317
rect 2385 6080 2390 6200
rect 2570 6080 2583 6200
rect 2385 6060 2583 6080
rect 2696 6020 2773 6215
rect 2805 8580 2882 8600
rect 2805 8460 2810 8580
rect 2870 8460 2882 8580
rect 2805 8445 2882 8460
rect 2995 8580 3193 8600
rect 2995 8460 3000 8580
rect 3180 8460 3193 8580
rect 2805 8343 2870 8445
rect 2805 6317 2882 8343
rect 2805 6215 2870 6317
rect 2805 6200 2882 6215
rect 2805 6080 2810 6200
rect 2870 6080 2882 6200
rect 2805 6060 2882 6080
rect 2995 6200 3193 8460
rect 3306 8445 3383 8640
rect 3319 8343 3383 8445
rect 3306 6317 3383 8343
rect 3318 6215 3383 6317
rect 2995 6080 3000 6200
rect 3180 6080 3193 6200
rect 2995 6060 3193 6080
rect 3306 6060 3383 6215
rect 3415 8445 3492 8640
rect 3605 8580 3803 8600
rect 3605 8460 3610 8580
rect 3790 8460 3803 8580
rect 3415 8343 3480 8445
rect 3415 6317 3492 8343
rect 3415 6215 3480 6317
rect 3415 6060 3492 6215
rect 3605 6200 3803 8460
rect 3916 8580 3993 8600
rect 3916 8460 3920 8580
rect 3980 8460 3993 8580
rect 3916 8445 3993 8460
rect 3929 8343 3993 8445
rect 3916 6317 3993 8343
rect 3928 6215 3993 6317
rect 3605 6080 3610 6200
rect 3790 6080 3803 6200
rect 3605 6060 3803 6080
rect 3916 6200 3993 6215
rect 3916 6080 3920 6200
rect 3980 6080 3993 6200
rect 3916 6060 3993 6080
rect 4025 8445 4102 8600
rect 4215 8580 4413 8600
rect 4215 8460 4220 8580
rect 4400 8460 4413 8580
rect 4025 8343 4090 8445
rect 4025 6317 4102 8343
rect 4025 6215 4090 6317
rect 2696 5900 2700 6020
rect 2760 5900 2773 6020
rect 2696 5880 2773 5900
rect 4025 6020 4102 6215
rect 4215 6200 4413 8460
rect 4526 8445 4603 8640
rect 4539 8343 4603 8445
rect 4526 6317 4603 8343
rect 4538 6215 4603 6317
rect 4215 6080 4220 6200
rect 4400 6080 4413 6200
rect 4215 6060 4413 6080
rect 4526 6060 4603 6215
rect 4635 8445 4712 8640
rect 4635 8343 4700 8445
rect 4635 6317 4712 8343
rect 4635 6215 4700 6317
rect 4025 5900 4030 6020
rect 4090 5900 4102 6020
rect 4025 5880 4102 5900
rect 4635 5840 4712 6215
rect 4825 5840 5023 8640
rect 5136 8445 5213 8640
rect 5149 8343 5213 8445
rect 5136 6317 5213 8343
rect 5148 6215 5213 6317
rect 5136 5840 5213 6215
rect 7690 8600 7770 8640
rect 7690 5880 7700 8600
rect 7760 5880 7770 8600
rect 7690 5840 7770 5880
rect 7815 8445 7892 8640
rect 7815 8343 7880 8445
rect 7815 6317 7892 8343
rect 7815 6215 7880 6317
rect 7815 5840 7892 6215
rect 8005 5840 8203 8640
rect 8316 8445 8393 8640
rect 8329 8343 8393 8445
rect 8316 6317 8393 8343
rect 8328 6215 8393 6317
rect 8316 5840 8393 6215
rect 8425 8445 8502 8640
rect 8615 8580 8813 8600
rect 8615 8460 8620 8580
rect 8800 8460 8813 8580
rect 8425 8343 8490 8445
rect 8425 6317 8502 8343
rect 8425 6215 8490 6317
rect 8425 6060 8502 6215
rect 8615 6200 8813 8460
rect 8926 8445 9003 8600
rect 8939 8343 9003 8445
rect 8926 6317 9003 8343
rect 8938 6215 9003 6317
rect 8615 6080 8620 6200
rect 8800 6080 8813 6200
rect 8615 6060 8813 6080
rect 8926 6020 9003 6215
rect 8926 5900 8930 6020
rect 8990 5900 9003 6020
rect 8926 5880 9003 5900
rect 9035 8445 9112 8600
rect 9225 8580 9423 8600
rect 9225 8460 9230 8580
rect 9410 8460 9423 8580
rect 9035 8343 9100 8445
rect 9035 6317 9112 8343
rect 9035 6215 9100 6317
rect 9035 6020 9112 6215
rect 9225 6200 9423 8460
rect 9536 8445 9613 8640
rect 9549 8343 9613 8445
rect 9536 6317 9613 8343
rect 9548 6215 9613 6317
rect 9225 6080 9230 6200
rect 9410 6080 9423 6200
rect 9225 6060 9423 6080
rect 9536 6060 9613 6215
rect 9645 8445 9722 8640
rect 9835 8580 10033 8600
rect 9835 8460 9840 8580
rect 10020 8460 10033 8580
rect 9645 8343 9710 8445
rect 9645 6317 9722 8343
rect 9645 6215 9710 6317
rect 9645 6060 9722 6215
rect 9835 6200 10033 8460
rect 10146 8445 10223 8600
rect 10159 8343 10223 8445
rect 10146 6317 10223 8343
rect 10158 6215 10223 6317
rect 9835 6080 9840 6200
rect 10020 6080 10033 6200
rect 9835 6060 10033 6080
rect 9035 5900 9040 6020
rect 9100 5900 9112 6020
rect 9035 5880 9112 5900
rect 10146 6020 10223 6215
rect 10146 5900 10150 6020
rect 10210 5900 10223 6020
rect 10146 5890 10223 5900
rect 10255 8445 10332 8600
rect 10445 8580 10643 8600
rect 10445 8460 10450 8580
rect 10630 8460 10643 8580
rect 10255 8343 10320 8445
rect 10255 6317 10332 8343
rect 10255 6215 10320 6317
rect 10255 6020 10332 6215
rect 10445 6200 10643 8460
rect 10756 8445 10833 8640
rect 10769 8343 10833 8445
rect 10756 6317 10833 8343
rect 10768 6215 10833 6317
rect 10445 6080 10450 6200
rect 10630 6080 10643 6200
rect 10445 6060 10643 6080
rect 10756 6060 10833 6215
rect 10865 8445 10942 8640
rect 11055 8580 11253 8600
rect 11055 8460 11060 8580
rect 11240 8460 11253 8580
rect 10865 8343 10930 8445
rect 10865 6317 10942 8343
rect 10865 6215 10930 6317
rect 10865 6060 10942 6215
rect 11055 6200 11253 8460
rect 11366 8445 11443 8600
rect 11379 8343 11443 8445
rect 11366 6317 11443 8343
rect 11378 6215 11443 6317
rect 11055 6080 11060 6200
rect 11240 6080 11253 6200
rect 11055 6060 11253 6080
rect 10255 5900 10260 6020
rect 10320 5900 10332 6020
rect 10255 5890 10332 5900
rect 11366 6020 11443 6215
rect 11475 8580 11552 8600
rect 11475 8460 11480 8580
rect 11540 8460 11552 8580
rect 11475 8445 11552 8460
rect 11665 8580 11863 8600
rect 11665 8460 11670 8580
rect 11850 8460 11863 8580
rect 11475 8343 11540 8445
rect 11475 6317 11552 8343
rect 11475 6215 11540 6317
rect 11475 6200 11552 6215
rect 11475 6080 11480 6200
rect 11540 6080 11552 6200
rect 11475 6060 11552 6080
rect 11665 6200 11863 8460
rect 11976 8445 12053 8640
rect 11989 8343 12053 8445
rect 11976 6317 12053 8343
rect 11988 6215 12053 6317
rect 11665 6080 11670 6200
rect 11850 6080 11863 6200
rect 11665 6060 11863 6080
rect 11976 6060 12053 6215
rect 12085 8445 12162 8640
rect 12275 8580 12473 8600
rect 12275 8460 12280 8580
rect 12460 8460 12473 8580
rect 12085 8343 12150 8445
rect 12085 6317 12162 8343
rect 12085 6215 12150 6317
rect 12085 6060 12162 6215
rect 12275 6200 12473 8460
rect 12586 8580 12663 8600
rect 12586 8460 12590 8580
rect 12650 8460 12663 8580
rect 12586 8445 12663 8460
rect 12599 8343 12663 8445
rect 12586 6317 12663 8343
rect 12598 6215 12663 6317
rect 12275 6080 12280 6200
rect 12460 6080 12473 6200
rect 12275 6060 12473 6080
rect 12586 6200 12663 6215
rect 12586 6080 12590 6200
rect 12650 6080 12663 6200
rect 12586 6060 12663 6080
rect 12695 8445 12772 8600
rect 12885 8580 13083 8600
rect 12885 8460 12890 8580
rect 13070 8460 13083 8580
rect 12695 8343 12760 8445
rect 12695 6317 12772 8343
rect 12695 6215 12760 6317
rect 11366 5900 11370 6020
rect 11430 5900 11443 6020
rect 11366 5890 11443 5900
rect 12695 6020 12772 6215
rect 12885 6200 13083 8460
rect 13196 8445 13273 8640
rect 13209 8343 13273 8445
rect 13196 6317 13273 8343
rect 13208 6215 13273 6317
rect 12885 6080 12890 6200
rect 13070 6080 13083 6200
rect 12885 6060 13083 6080
rect 13196 6060 13273 6215
rect 13305 8445 13382 8640
rect 13495 8580 13693 8600
rect 13495 8460 13500 8580
rect 13680 8460 13693 8580
rect 13305 8343 13370 8445
rect 13305 6317 13382 8343
rect 13305 6215 13370 6317
rect 13305 6060 13382 6215
rect 13495 6200 13693 8460
rect 13806 8445 13883 8600
rect 13819 8343 13883 8445
rect 13806 6317 13883 8343
rect 13818 6215 13883 6317
rect 13495 6080 13500 6200
rect 13680 6080 13693 6200
rect 13495 6060 13693 6080
rect 12695 5900 12700 6020
rect 12760 5900 12772 6020
rect 12695 5890 12772 5900
rect 13806 6020 13883 6215
rect 13806 5900 13810 6020
rect 13870 5900 13883 6020
rect 13806 5890 13883 5900
rect 13915 8445 13992 8600
rect 14105 8580 14303 8600
rect 14105 8460 14110 8580
rect 14290 8460 14303 8580
rect 13915 8343 13980 8445
rect 13915 6317 13992 8343
rect 13915 6215 13980 6317
rect 13915 6020 13992 6215
rect 13915 5900 13920 6020
rect 13980 5900 13992 6020
rect 13915 5890 13992 5900
rect 14105 6200 14303 8460
rect 14416 8445 14493 8640
rect 14429 8343 14493 8445
rect 14416 6317 14493 8343
rect 14428 6215 14493 6317
rect 14105 6080 14110 6200
rect 14290 6080 14303 6200
rect 14105 5890 14303 6080
rect 14416 6060 14493 6215
rect 14525 8445 14602 8640
rect 14715 8580 14913 8600
rect 14715 8460 14720 8580
rect 14900 8460 14913 8580
rect 14525 8343 14590 8445
rect 14525 6317 14602 8343
rect 14525 6215 14590 6317
rect 14525 6060 14602 6215
rect 14715 6200 14913 8460
rect 15026 8445 15103 8600
rect 15039 8343 15103 8445
rect 15026 6317 15103 8343
rect 15038 6215 15103 6317
rect 14715 6080 14720 6200
rect 14900 6080 14913 6200
rect 14715 6060 14913 6080
rect 15026 6020 15103 6215
rect 15026 5900 15030 6020
rect 15090 5900 15103 6020
rect 15026 5890 15103 5900
rect 15135 8445 15212 8600
rect 15325 8580 15523 8600
rect 15325 8460 15330 8580
rect 15510 8460 15523 8580
rect 15135 8343 15200 8445
rect 15135 6317 15212 8343
rect 15135 6215 15200 6317
rect 15135 6020 15212 6215
rect 15325 6200 15523 8460
rect 15636 8445 15713 8640
rect 15649 8343 15713 8445
rect 15636 6317 15713 8343
rect 15648 6215 15713 6317
rect 15325 6080 15330 6200
rect 15510 6080 15523 6200
rect 15325 6060 15523 6080
rect 15636 6060 15713 6215
rect 15745 8445 15822 8640
rect 15745 8343 15810 8445
rect 15745 6317 15822 8343
rect 15745 6215 15810 6317
rect 15135 5900 15140 6020
rect 15200 5900 15212 6020
rect 15135 5890 15212 5900
rect 15745 5840 15822 6215
rect 15935 5840 16133 8640
rect 16246 8600 16500 8640
rect 16246 8445 16370 8600
rect 16259 8343 16370 8445
rect 16246 6317 16370 8343
rect 16258 6215 16370 6317
rect 16246 5880 16370 6215
rect 16420 5880 16500 8600
rect 16246 5840 16500 5880
rect -1490 5830 16500 5840
rect -1490 5780 -860 5830
rect 7650 5780 7810 5830
rect 16320 5780 16500 5830
rect -1490 5570 16500 5780
rect -1490 5490 10040 5570
rect 15450 5490 16500 5570
rect -1490 5450 16500 5490
rect 9390 5370 16500 5450
rect 170 4990 8830 5350
rect 170 4940 1120 4990
rect 8350 4940 8830 4990
rect -1490 4500 90 4510
rect -1490 4380 -230 4500
rect 80 4380 90 4500
rect -1490 4370 90 4380
rect -1490 3810 -990 4370
rect -1490 140 -990 700
rect -1490 130 90 140
rect -1490 10 -230 130
rect 80 10 90 130
rect -1490 0 90 10
rect 170 -370 440 4940
rect 590 4930 8830 4940
rect 590 4880 1660 4930
rect 7810 4883 8830 4930
rect 590 -370 970 4880
rect 1020 4870 1660 4880
rect 1020 4365 1172 4870
rect 1020 4258 1153 4365
rect 1020 258 1172 4258
rect 1020 151 1153 258
rect 1020 -340 1172 151
rect 1265 -340 1491 4870
rect 1584 4365 1660 4870
rect 1603 4258 1660 4365
rect 1584 258 1660 4258
rect 1603 151 1660 258
rect 1584 -340 1660 151
rect 1020 -370 1660 -340
rect 1706 4680 1782 4883
rect 1706 4560 1710 4680
rect 1780 4560 1782 4680
rect 1706 4365 1782 4560
rect 1706 4258 1763 4365
rect 1706 258 1782 4258
rect 1706 151 1763 258
rect 1706 -368 1782 151
rect 1875 130 2101 4883
rect 2194 4365 2270 4883
rect 2213 4258 2270 4365
rect 2194 258 2270 4258
rect 2213 151 2270 258
rect 1875 10 1880 130
rect 2090 10 2101 130
rect 1875 -368 2101 10
rect 2194 -50 2270 151
rect 2194 -170 2200 -50
rect 2194 -368 2270 -170
rect 2316 4680 2392 4883
rect 2316 4560 2320 4680
rect 2390 4560 2392 4680
rect 2316 4365 2392 4560
rect 2316 4258 2373 4365
rect 2316 258 2392 4258
rect 2316 151 2373 258
rect 2316 -368 2392 151
rect 2485 130 2711 4883
rect 2804 4365 2880 4883
rect 2823 4258 2880 4365
rect 2804 258 2880 4258
rect 2823 151 2880 258
rect 2485 10 2490 130
rect 2700 10 2711 130
rect 2485 -368 2711 10
rect 2804 -50 2880 151
rect 2804 -170 2810 -50
rect 2804 -368 2880 -170
rect 2926 4860 3002 4883
rect 2926 4740 2930 4860
rect 3000 4740 3002 4860
rect 2926 4365 3002 4740
rect 3095 4500 3321 4883
rect 3095 4380 3100 4500
rect 3310 4380 3321 4500
rect 2926 4258 2983 4365
rect 2926 258 3002 4258
rect 2926 151 2983 258
rect 2926 -368 3002 151
rect 3095 -368 3321 4380
rect 3414 4365 3490 4883
rect 3433 4258 3490 4365
rect 3414 258 3490 4258
rect 3433 151 3490 258
rect 3414 -230 3490 151
rect 3414 -350 3420 -230
rect 3414 -368 3490 -350
rect 3536 4365 3612 4883
rect 3536 4258 3593 4365
rect 3536 258 3612 4258
rect 3536 151 3593 258
rect 3536 -50 3612 151
rect 3536 -170 3540 -50
rect 3610 -170 3612 -50
rect 3536 -368 3612 -170
rect 3705 130 3931 4883
rect 4024 4680 4100 4883
rect 4024 4560 4030 4680
rect 4024 4365 4100 4560
rect 4043 4258 4100 4365
rect 4024 258 4100 4258
rect 4043 151 4100 258
rect 3705 10 3710 130
rect 3920 10 3931 130
rect 3705 -368 3931 10
rect 4024 -368 4100 151
rect 4146 4365 4222 4883
rect 4315 4500 4541 4883
rect 4315 4380 4320 4500
rect 4530 4380 4541 4500
rect 4146 4258 4203 4365
rect 4146 258 4222 4258
rect 4146 151 4203 258
rect 4146 -230 4222 151
rect 4146 -350 4150 -230
rect 4220 -350 4222 -230
rect 4146 -368 4222 -350
rect 4315 -368 4541 4380
rect 4634 4860 4710 4883
rect 4634 4740 4640 4860
rect 4634 4365 4710 4740
rect 4653 4258 4710 4365
rect 4634 258 4710 4258
rect 4653 151 4710 258
rect 4634 -368 4710 151
rect 4756 4860 4832 4883
rect 4756 4740 4760 4860
rect 4830 4740 4832 4860
rect 4756 4365 4832 4740
rect 4925 4500 5151 4883
rect 4925 4380 4930 4500
rect 5140 4380 5151 4500
rect 4756 4258 4813 4365
rect 4756 258 4832 4258
rect 4756 151 4813 258
rect 4756 -368 4832 151
rect 4925 -368 5151 4380
rect 5244 4365 5320 4883
rect 5263 4258 5320 4365
rect 5244 258 5320 4258
rect 5263 151 5320 258
rect 5244 -230 5320 151
rect 5244 -350 5250 -230
rect 5244 -368 5320 -350
rect 5366 4680 5442 4883
rect 5366 4560 5370 4680
rect 5440 4560 5442 4680
rect 5366 4365 5442 4560
rect 5366 4258 5423 4365
rect 5366 258 5442 4258
rect 5366 151 5423 258
rect 5366 -368 5442 151
rect 5535 130 5761 4883
rect 5854 4365 5930 4883
rect 5873 4258 5930 4365
rect 5854 258 5930 4258
rect 5873 151 5930 258
rect 5535 10 5540 130
rect 5750 10 5761 130
rect 5535 -368 5761 10
rect 5854 -50 5930 151
rect 5854 -170 5860 -50
rect 5854 -368 5930 -170
rect 5976 4365 6052 4883
rect 6145 4500 6371 4883
rect 6145 4380 6150 4500
rect 6360 4380 6371 4500
rect 5976 4258 6033 4365
rect 5976 258 6052 4258
rect 5976 151 6033 258
rect 5976 -230 6052 151
rect 5976 -350 5980 -230
rect 6050 -350 6052 -230
rect 5976 -368 6052 -350
rect 6145 -368 6371 4380
rect 6464 4860 6540 4883
rect 6464 4740 6470 4860
rect 6464 4365 6540 4740
rect 6483 4258 6540 4365
rect 6464 258 6540 4258
rect 6483 151 6540 258
rect 6464 -368 6540 151
rect 6586 4365 6662 4883
rect 6586 4258 6643 4365
rect 6586 258 6662 4258
rect 6586 151 6643 258
rect 6586 -50 6662 151
rect 6586 -170 6590 -50
rect 6660 -170 6662 -50
rect 6586 -368 6662 -170
rect 6755 130 6981 4883
rect 7074 4680 7150 4883
rect 7074 4560 7080 4680
rect 7074 4365 7150 4560
rect 7093 4258 7150 4365
rect 7074 258 7150 4258
rect 7093 151 7150 258
rect 6755 10 6760 130
rect 6970 10 6981 130
rect 6755 -368 6981 10
rect 7074 -368 7150 151
rect 7196 4365 7272 4883
rect 7365 4500 7591 4883
rect 7365 4380 7370 4500
rect 7580 4380 7591 4500
rect 7196 4258 7253 4365
rect 7196 258 7272 4258
rect 7196 151 7253 258
rect 7196 -230 7272 151
rect 7196 -350 7200 -230
rect 7270 -350 7272 -230
rect 7196 -368 7272 -350
rect 7365 -368 7591 4380
rect 7684 4860 7760 4883
rect 7684 4740 7690 4860
rect 7684 4365 7760 4740
rect 7703 4258 7760 4365
rect 7684 258 7760 4258
rect 7703 151 7760 258
rect 7684 -368 7760 151
rect 7806 4880 8830 4883
rect 7806 4870 8450 4880
rect 7806 4365 7882 4870
rect 7806 4258 7863 4365
rect 7806 258 7882 4258
rect 7806 151 7863 258
rect 7806 -350 7882 151
rect 7975 -350 8201 4870
rect 8294 4365 8450 4870
rect 8313 4258 8450 4365
rect 8294 258 8450 4258
rect 8313 151 8450 258
rect 8294 -350 8450 151
rect 7806 -368 8450 -350
rect -1490 -410 1660 -370
rect 7810 -370 8450 -368
rect 8500 -370 8830 4880
rect 9390 5320 9770 5370
rect 15970 5320 16500 5370
rect 9390 5270 16500 5320
rect 9390 340 9670 5270
rect 9720 5130 16020 5270
rect 9720 4800 9850 5130
rect 10310 5070 10470 5130
rect 10930 5070 11090 5130
rect 11550 5070 11710 5130
rect 12170 5070 12330 5130
rect 12790 5070 12950 5130
rect 13410 5070 13570 5130
rect 14030 5070 14190 5130
rect 14650 5070 14810 5130
rect 15270 5070 15430 5130
rect 15890 5070 16020 5130
rect 9878 5050 9970 5060
rect 9878 4930 9880 5050
rect 9960 4930 9970 5050
rect 9878 4828 9970 4930
rect 9720 800 9868 4800
rect 9720 530 9850 800
rect 9896 772 9952 4828
rect 9998 4800 10160 5070
rect 10188 5050 10280 5070
rect 10188 4930 10190 5050
rect 10270 4930 10280 5050
rect 10188 4828 10280 4930
rect 9980 800 10178 4800
rect 9878 670 9970 772
rect 9878 550 9880 670
rect 9960 550 9970 670
rect 9878 530 9970 550
rect 9720 340 9800 530
rect 9998 490 10160 800
rect 10206 772 10262 4828
rect 10308 4800 10470 5070
rect 10498 5050 10590 5070
rect 10498 4930 10500 5050
rect 10580 4930 10590 5050
rect 10498 4828 10590 4930
rect 10290 800 10488 4800
rect 10188 670 10280 772
rect 10188 550 10190 670
rect 10270 550 10280 670
rect 10188 530 10280 550
rect 10308 530 10470 800
rect 10516 772 10572 4828
rect 10618 4800 10780 5070
rect 10808 5050 10900 5070
rect 10808 4930 10810 5050
rect 10890 4930 10900 5050
rect 10808 4828 10900 4930
rect 10600 800 10798 4800
rect 10498 670 10590 772
rect 10498 550 10500 670
rect 10580 550 10590 670
rect 10498 530 10590 550
rect 9998 370 10010 490
rect 10150 370 10160 490
rect 9998 350 10160 370
rect 10618 490 10780 800
rect 10826 772 10882 4828
rect 10928 4800 11090 5070
rect 11118 5050 11210 5070
rect 11118 4930 11120 5050
rect 11200 4930 11210 5050
rect 11118 4828 11210 4930
rect 10910 800 11108 4800
rect 10808 670 10900 772
rect 10808 550 10810 670
rect 10890 550 10900 670
rect 10808 530 10900 550
rect 10928 530 11090 800
rect 11136 772 11192 4828
rect 11238 4800 11400 5070
rect 11428 5050 11520 5070
rect 11428 4930 11430 5050
rect 11510 4930 11520 5050
rect 11428 4828 11520 4930
rect 11220 800 11418 4800
rect 11118 670 11210 772
rect 11118 550 11120 670
rect 11200 550 11210 670
rect 11118 530 11210 550
rect 10618 370 10630 490
rect 10770 370 10780 490
rect 10618 350 10780 370
rect 11238 490 11400 800
rect 11446 772 11502 4828
rect 11548 4800 11710 5070
rect 11738 5050 11830 5070
rect 11738 4930 11740 5050
rect 11820 4930 11830 5050
rect 11738 4828 11830 4930
rect 11530 800 11728 4800
rect 11428 670 11520 772
rect 11428 550 11430 670
rect 11510 550 11520 670
rect 11428 530 11520 550
rect 11548 530 11710 800
rect 11756 772 11812 4828
rect 11858 4800 12020 5070
rect 12048 5050 12140 5070
rect 12048 4930 12050 5050
rect 12130 4930 12140 5050
rect 12048 4828 12140 4930
rect 11840 800 12038 4800
rect 11738 670 11830 772
rect 11738 550 11740 670
rect 11820 550 11830 670
rect 11738 530 11830 550
rect 11238 370 11250 490
rect 11390 370 11400 490
rect 11238 350 11400 370
rect 11858 490 12020 800
rect 12066 772 12122 4828
rect 12168 4800 12330 5070
rect 12358 5050 12450 5070
rect 12358 4930 12360 5050
rect 12440 4930 12450 5050
rect 12358 4828 12450 4930
rect 12150 800 12348 4800
rect 12048 670 12140 772
rect 12048 550 12050 670
rect 12130 550 12140 670
rect 12048 530 12140 550
rect 12168 530 12330 800
rect 12376 772 12432 4828
rect 12478 4800 12640 5070
rect 12668 5050 12760 5070
rect 12668 4930 12670 5050
rect 12750 4930 12760 5050
rect 12668 4828 12760 4930
rect 12460 800 12658 4800
rect 12358 670 12450 772
rect 12358 550 12360 670
rect 12440 550 12450 670
rect 12358 530 12450 550
rect 11858 370 11870 490
rect 12010 370 12020 490
rect 11858 350 12020 370
rect 12478 490 12640 800
rect 12686 772 12742 4828
rect 12788 4800 12950 5070
rect 12978 5050 13070 5070
rect 12978 4930 12980 5050
rect 13060 4930 13070 5050
rect 12978 4828 13070 4930
rect 12770 800 12968 4800
rect 12668 670 12760 772
rect 12668 550 12670 670
rect 12750 550 12760 670
rect 12668 530 12760 550
rect 12788 530 12950 800
rect 12996 772 13052 4828
rect 13098 4800 13260 5070
rect 13288 5050 13380 5070
rect 13288 4930 13290 5050
rect 13370 4930 13380 5050
rect 13288 4828 13380 4930
rect 13080 800 13278 4800
rect 12978 670 13070 772
rect 12978 550 12980 670
rect 13060 550 13070 670
rect 12978 530 13070 550
rect 12478 370 12490 490
rect 12630 370 12640 490
rect 12478 350 12640 370
rect 13098 490 13260 800
rect 13306 772 13362 4828
rect 13408 4800 13570 5070
rect 13598 5050 13690 5070
rect 13598 4930 13600 5050
rect 13680 4930 13690 5050
rect 13598 4828 13690 4930
rect 13390 800 13588 4800
rect 13288 670 13380 772
rect 13288 550 13290 670
rect 13370 550 13380 670
rect 13288 530 13380 550
rect 13408 530 13570 800
rect 13616 772 13672 4828
rect 13718 4800 13880 5070
rect 13908 5050 14000 5070
rect 13908 4930 13910 5050
rect 13990 4930 14000 5050
rect 13908 4828 14000 4930
rect 13700 800 13898 4800
rect 13598 670 13690 772
rect 13598 550 13600 670
rect 13680 550 13690 670
rect 13598 530 13690 550
rect 13098 370 13110 490
rect 13250 370 13260 490
rect 13098 350 13260 370
rect 13718 490 13880 800
rect 13926 772 13982 4828
rect 14028 4800 14190 5070
rect 14218 5050 14310 5070
rect 14218 4930 14220 5050
rect 14300 4930 14310 5050
rect 14218 4828 14310 4930
rect 14010 800 14208 4800
rect 13908 670 14000 772
rect 13908 550 13910 670
rect 13990 550 14000 670
rect 13908 530 14000 550
rect 14028 530 14190 800
rect 14236 772 14292 4828
rect 14338 4800 14500 5070
rect 14528 5050 14620 5070
rect 14528 4930 14530 5050
rect 14610 4930 14620 5050
rect 14528 4828 14620 4930
rect 14320 800 14518 4800
rect 14218 670 14310 772
rect 14218 550 14220 670
rect 14300 550 14310 670
rect 14218 530 14310 550
rect 13718 370 13730 490
rect 13870 370 13880 490
rect 13718 350 13880 370
rect 14338 490 14500 800
rect 14546 772 14602 4828
rect 14648 4800 14810 5070
rect 14838 5050 14930 5070
rect 14838 4930 14840 5050
rect 14920 4930 14930 5050
rect 14838 4828 14930 4930
rect 14630 800 14828 4800
rect 14528 670 14620 772
rect 14528 550 14530 670
rect 14610 550 14620 670
rect 14528 530 14620 550
rect 14648 530 14810 800
rect 14856 772 14912 4828
rect 14958 4800 15120 5070
rect 15148 5050 15240 5070
rect 15148 4930 15150 5050
rect 15230 4930 15240 5050
rect 15148 4828 15240 4930
rect 14940 800 15138 4800
rect 14838 670 14930 772
rect 14838 550 14840 670
rect 14920 550 14930 670
rect 14838 530 14930 550
rect 14338 370 14350 490
rect 14490 370 14500 490
rect 14338 350 14500 370
rect 14958 490 15120 800
rect 15166 772 15222 4828
rect 15268 4800 15430 5070
rect 15458 5050 15550 5070
rect 15458 4930 15460 5050
rect 15540 4930 15550 5050
rect 15458 4828 15550 4930
rect 15250 800 15448 4800
rect 15148 670 15240 772
rect 15148 550 15150 670
rect 15230 550 15240 670
rect 15148 530 15240 550
rect 15268 530 15430 800
rect 15476 772 15532 4828
rect 15578 4800 15740 5070
rect 15768 5050 15860 5060
rect 15768 4930 15770 5050
rect 15850 4930 15860 5050
rect 15768 4828 15860 4930
rect 15560 800 15758 4800
rect 15458 670 15550 772
rect 15458 550 15460 670
rect 15540 550 15550 670
rect 15458 530 15550 550
rect 14958 370 14970 490
rect 15110 370 15120 490
rect 14958 350 15120 370
rect 15578 490 15740 800
rect 15786 772 15842 4828
rect 15888 4800 16020 5070
rect 15870 800 16020 4800
rect 15768 670 15860 772
rect 15768 550 15770 670
rect 15850 550 15860 670
rect 15768 530 15860 550
rect 15888 530 16020 800
rect 15578 370 15590 490
rect 15730 370 15740 490
rect 15578 350 15740 370
rect 9390 300 9800 340
rect 15930 340 16020 530
rect 16070 5130 16500 5270
rect 16070 340 16410 5130
rect 15930 300 16410 340
rect 9390 290 16410 300
rect 9390 240 9770 290
rect 15970 240 16410 290
rect 9390 -40 16410 240
rect 16690 820 17520 830
rect 16690 350 16700 820
rect 17510 350 17520 820
rect 16690 -270 17520 350
rect 7810 -410 8830 -370
rect -1490 -420 8830 -410
rect -1490 -470 1120 -420
rect 8350 -470 8830 -420
rect -1490 -780 8830 -470
rect 9060 -280 17520 -270
rect 9060 -580 9070 -280
rect 9590 -580 17520 -280
rect 9060 -590 17520 -580
rect -1490 -1650 590 -780
rect 11430 -800 14960 -790
rect 11430 -1010 11440 -800
rect 11840 -1010 12050 -800
rect 12450 -1010 12670 -800
rect 13070 -1010 13300 -800
rect 13690 -1010 14960 -800
rect 11430 -1020 14960 -1010
rect 14310 -1148 14490 -1080
rect 6090 -1170 8300 -1160
rect 6090 -1550 6100 -1170
rect 6640 -1550 7730 -1170
rect 8270 -1550 8300 -1170
rect 6090 -1560 8300 -1550
rect 14310 -1498 14416 -1148
rect 14450 -1498 14490 -1148
rect 14560 -1450 14960 -1020
rect 15351 -1030 17520 -790
rect 15351 -1454 15772 -1030
rect 15860 -1148 16050 -1080
rect 14310 -1550 14490 -1498
rect 15860 -1498 15874 -1148
rect 15908 -1498 16050 -1148
rect 15860 -1550 16050 -1498
rect 14310 -1560 16050 -1550
rect 8440 -1594 14512 -1560
rect 15812 -1594 16510 -1560
rect 8440 -1650 16510 -1594
rect -1490 -1770 16510 -1650
rect -1490 -1820 7760 -1770
rect 16330 -1820 16510 -1770
rect -1490 -1830 16510 -1820
rect -1490 -1870 7720 -1830
rect -1490 -1950 7660 -1870
rect -1490 -2000 -1160 -1950
rect 7410 -2000 7660 -1950
rect -1490 -2010 7660 -2000
rect -1490 -2050 -1054 -2010
rect -1490 -4790 -1260 -2050
rect -1210 -2406 -1054 -2050
rect -1210 -2508 -1066 -2406
rect -1210 -4516 -1054 -2508
rect -1210 -4618 -1066 -4516
rect -1210 -4790 -1054 -4618
rect -1490 -4830 -1054 -4790
rect -936 -4830 -748 -2010
rect -630 -2406 -553 -2010
rect -20 -2090 57 -2070
rect 50 -2210 57 -2090
rect -618 -2508 -553 -2406
rect -630 -4516 -553 -2508
rect -618 -4618 -553 -4516
rect -630 -4830 -553 -4618
rect -521 -2406 -444 -2250
rect -326 -2270 -138 -2250
rect -326 -2390 -320 -2270
rect -150 -2390 -138 -2270
rect -521 -2508 -456 -2406
rect -521 -4516 -444 -2508
rect -521 -4618 -456 -4516
rect -521 -4830 -444 -4618
rect -326 -4630 -138 -2390
rect -20 -2406 57 -2210
rect -8 -2508 57 -2406
rect -20 -4516 57 -2508
rect -8 -4618 57 -4516
rect -326 -4750 -320 -4630
rect -150 -4750 -138 -4630
rect -326 -4770 -138 -4750
rect -20 -4770 57 -4618
rect 89 -2090 166 -2070
rect 89 -2210 90 -2090
rect 160 -2210 166 -2090
rect 89 -2406 166 -2210
rect 1200 -2090 1277 -2070
rect 1270 -2210 1277 -2090
rect 284 -2270 472 -2250
rect 284 -2390 290 -2270
rect 460 -2390 472 -2270
rect 89 -2508 154 -2406
rect 89 -4516 166 -2508
rect 89 -4618 154 -4516
rect 89 -4770 166 -4618
rect 284 -4630 472 -2390
rect 590 -2406 667 -2250
rect 602 -2508 667 -2406
rect 590 -4516 667 -2508
rect 602 -4618 667 -4516
rect 284 -4750 290 -4630
rect 460 -4750 472 -4630
rect 284 -4770 472 -4750
rect 590 -4830 667 -4618
rect 699 -2406 776 -2250
rect 894 -2270 1082 -2250
rect 894 -2390 900 -2270
rect 1070 -2390 1082 -2270
rect 699 -2508 764 -2406
rect 699 -4516 776 -2508
rect 699 -4618 764 -4516
rect 699 -4830 776 -4618
rect 894 -4630 1082 -2390
rect 1200 -2406 1277 -2210
rect 1212 -2508 1277 -2406
rect 1200 -4516 1277 -2508
rect 1212 -4618 1277 -4516
rect 894 -4750 900 -4630
rect 1070 -4750 1082 -4630
rect 894 -4770 1082 -4750
rect 1200 -4770 1277 -4618
rect 1309 -2090 1386 -2070
rect 1309 -2210 1310 -2090
rect 1380 -2210 1386 -2090
rect 1309 -2406 1386 -2210
rect 2420 -2090 2497 -2070
rect 2490 -2210 2497 -2090
rect 1504 -2270 1692 -2250
rect 1504 -2390 1510 -2270
rect 1680 -2390 1692 -2270
rect 1309 -2508 1374 -2406
rect 1309 -4516 1386 -2508
rect 1309 -4618 1374 -4516
rect 1309 -4770 1386 -4618
rect 1504 -4630 1692 -2390
rect 1810 -2406 1887 -2250
rect 1822 -2508 1887 -2406
rect 1810 -4516 1887 -2508
rect 1822 -4618 1887 -4516
rect 1504 -4750 1510 -4630
rect 1680 -4750 1692 -4630
rect 1504 -4770 1692 -4750
rect 1810 -4830 1887 -4618
rect 1919 -2406 1996 -2250
rect 2114 -2270 2302 -2250
rect 2114 -2390 2120 -2270
rect 2290 -2390 2302 -2270
rect 1919 -2508 1984 -2406
rect 1919 -4516 1996 -2508
rect 1919 -4618 1984 -4516
rect 1919 -4830 1996 -4618
rect 2114 -4630 2302 -2390
rect 2420 -2406 2497 -2210
rect 3749 -2090 3826 -2070
rect 3749 -2210 3750 -2090
rect 3820 -2210 3826 -2090
rect 2432 -2508 2497 -2406
rect 2420 -4516 2497 -2508
rect 2432 -4618 2497 -4516
rect 2114 -4750 2120 -4630
rect 2290 -4750 2302 -4630
rect 2114 -4770 2302 -4750
rect 2420 -4770 2497 -4618
rect 2529 -2270 2606 -2250
rect 2529 -2390 2530 -2270
rect 2600 -2390 2606 -2270
rect 2529 -2406 2606 -2390
rect 2724 -2270 2912 -2250
rect 2724 -2390 2730 -2270
rect 2900 -2390 2912 -2270
rect 2529 -2508 2594 -2406
rect 2529 -4516 2606 -2508
rect 2529 -4618 2594 -4516
rect 2529 -4630 2606 -4618
rect 2529 -4750 2530 -4630
rect 2600 -4750 2606 -4630
rect 2529 -4770 2606 -4750
rect 2724 -4630 2912 -2390
rect 3030 -2406 3107 -2250
rect 3042 -2508 3107 -2406
rect 3030 -4516 3107 -2508
rect 3042 -4618 3107 -4516
rect 2724 -4750 2730 -4630
rect 2900 -4750 2912 -4630
rect 2724 -4770 2912 -4750
rect 3030 -4830 3107 -4618
rect 3139 -2406 3216 -2250
rect 3334 -2270 3522 -2250
rect 3334 -2390 3340 -2270
rect 3510 -2390 3522 -2270
rect 3139 -2508 3204 -2406
rect 3139 -4516 3216 -2508
rect 3139 -4618 3204 -4516
rect 3139 -4830 3216 -4618
rect 3334 -4630 3522 -2390
rect 3640 -2270 3717 -2250
rect 3710 -2390 3717 -2270
rect 3640 -2406 3717 -2390
rect 3652 -2508 3717 -2406
rect 3640 -4516 3717 -2508
rect 3652 -4618 3717 -4516
rect 3334 -4750 3340 -4630
rect 3510 -4750 3522 -4630
rect 3334 -4770 3522 -4750
rect 3640 -4630 3717 -4618
rect 3710 -4750 3717 -4630
rect 3640 -4770 3717 -4750
rect 3749 -2406 3826 -2210
rect 4860 -2090 4937 -2070
rect 4930 -2210 4937 -2090
rect 3944 -2270 4132 -2250
rect 3944 -2390 3950 -2270
rect 4120 -2390 4132 -2270
rect 3749 -2508 3814 -2406
rect 3749 -4516 3826 -2508
rect 3749 -4618 3814 -4516
rect 3749 -4770 3826 -4618
rect 3944 -4630 4132 -2390
rect 4250 -2406 4327 -2250
rect 4262 -2508 4327 -2406
rect 4250 -4516 4327 -2508
rect 4262 -4618 4327 -4516
rect 3944 -4750 3950 -4630
rect 4120 -4750 4132 -4630
rect 3944 -4770 4132 -4750
rect 4250 -4830 4327 -4618
rect 4359 -2406 4436 -2250
rect 4554 -2270 4742 -2250
rect 4554 -2390 4560 -2270
rect 4730 -2390 4742 -2270
rect 4359 -2508 4424 -2406
rect 4359 -4516 4436 -2508
rect 4359 -4618 4424 -4516
rect 4359 -4830 4436 -4618
rect 4554 -4630 4742 -2390
rect 4860 -2406 4937 -2210
rect 4872 -2508 4937 -2406
rect 4860 -4516 4937 -2508
rect 4872 -4618 4937 -4516
rect 4554 -4750 4560 -4630
rect 4730 -4750 4742 -4630
rect 4554 -4770 4742 -4750
rect 4860 -4770 4937 -4618
rect 4969 -2090 5046 -2070
rect 4969 -2210 4970 -2090
rect 5040 -2210 5046 -2090
rect 4969 -2406 5046 -2210
rect 6080 -2090 6157 -2070
rect 6150 -2210 6157 -2090
rect 5164 -2270 5352 -2250
rect 5164 -2390 5170 -2270
rect 5340 -2390 5352 -2270
rect 4969 -2508 5034 -2406
rect 4969 -4516 5046 -2508
rect 4969 -4618 5034 -4516
rect 4969 -4770 5046 -4618
rect 5164 -4630 5352 -2390
rect 5470 -2406 5547 -2250
rect 5482 -2508 5547 -2406
rect 5470 -4516 5547 -2508
rect 5482 -4618 5547 -4516
rect 5164 -4750 5170 -4630
rect 5340 -4750 5352 -4630
rect 5164 -4770 5352 -4750
rect 5470 -4830 5547 -4618
rect 5579 -2406 5656 -2250
rect 5774 -2270 5962 -2250
rect 5774 -2390 5780 -2270
rect 5950 -2390 5962 -2270
rect 5579 -2508 5644 -2406
rect 5579 -4516 5656 -2508
rect 5579 -4618 5644 -4516
rect 5579 -4830 5656 -4618
rect 5774 -4630 5962 -2390
rect 6080 -2406 6157 -2210
rect 6092 -2508 6157 -2406
rect 6080 -4516 6157 -2508
rect 6092 -4618 6157 -4516
rect 5774 -4750 5780 -4630
rect 5950 -4750 5962 -4630
rect 5774 -4770 5962 -4750
rect 6080 -4770 6157 -4618
rect 6189 -2090 6266 -2070
rect 6189 -2210 6190 -2090
rect 6260 -2210 6266 -2090
rect 6189 -2406 6266 -2210
rect 6384 -2270 6572 -2250
rect 6384 -2390 6390 -2270
rect 6560 -2390 6572 -2270
rect 6189 -2508 6254 -2406
rect 6189 -4516 6266 -2508
rect 6189 -4618 6254 -4516
rect 6189 -4770 6266 -4618
rect 6384 -4630 6572 -2390
rect 6690 -2406 6767 -2250
rect 6702 -2508 6767 -2406
rect 6690 -4516 6767 -2508
rect 6702 -4618 6767 -4516
rect 6384 -4750 6390 -4630
rect 6560 -4750 6572 -4630
rect 6384 -4770 6572 -4750
rect 6690 -4830 6767 -4618
rect 6799 -2406 6876 -2010
rect 6799 -2508 6864 -2406
rect 6799 -4516 6876 -2508
rect 6799 -4618 6864 -4516
rect 6799 -4830 6876 -4618
rect 6994 -4830 7182 -2010
rect 7300 -2406 7377 -2010
rect 7312 -2508 7377 -2406
rect 7300 -4516 7377 -2508
rect 7312 -4618 7377 -4516
rect 7300 -4830 7377 -4618
rect 7450 -2050 7660 -2010
rect 7450 -4790 7460 -2050
rect 7510 -4790 7660 -2050
rect 7710 -4790 7720 -1870
rect 7450 -4830 7720 -4790
rect 7789 -2406 7866 -1830
rect 7789 -2508 7854 -2406
rect 7789 -4516 7866 -2508
rect 7789 -4618 7854 -4516
rect 7789 -4830 7866 -4618
rect 7984 -4830 8172 -1830
rect 8290 -2406 8367 -1830
rect 8900 -1910 8977 -1890
rect 8970 -2030 8977 -1910
rect 8302 -2508 8367 -2406
rect 8290 -4516 8367 -2508
rect 8302 -4618 8367 -4516
rect 8290 -4830 8367 -4618
rect 8399 -2406 8476 -2250
rect 8594 -2270 8782 -2250
rect 8594 -2390 8600 -2270
rect 8770 -2390 8782 -2270
rect 8399 -2508 8464 -2406
rect 8399 -4516 8476 -2508
rect 8399 -4618 8464 -4516
rect 8399 -4830 8476 -4618
rect 8594 -4630 8782 -2390
rect 8900 -2406 8977 -2030
rect 8912 -2508 8977 -2406
rect 8900 -4516 8977 -2508
rect 8912 -4618 8977 -4516
rect 8594 -4750 8600 -4630
rect 8770 -4750 8782 -4630
rect 8594 -4770 8782 -4750
rect 8900 -4770 8977 -4618
rect 9009 -1910 9086 -1890
rect 9009 -2030 9010 -1910
rect 9080 -2030 9086 -1910
rect 9009 -2406 9086 -2030
rect 10120 -1910 10197 -1890
rect 10190 -2030 10197 -1910
rect 9204 -2270 9392 -2250
rect 9204 -2390 9210 -2270
rect 9380 -2390 9392 -2270
rect 9009 -2508 9074 -2406
rect 9009 -4516 9086 -2508
rect 9009 -4618 9074 -4516
rect 9009 -4770 9086 -4618
rect 9204 -4630 9392 -2390
rect 9510 -2406 9587 -2250
rect 9522 -2508 9587 -2406
rect 9510 -4516 9587 -2508
rect 9522 -4618 9587 -4516
rect 9204 -4750 9210 -4630
rect 9380 -4750 9392 -4630
rect 9204 -4770 9392 -4750
rect 9510 -4830 9587 -4618
rect 9619 -2406 9696 -2250
rect 9814 -2270 10002 -2250
rect 9814 -2390 9820 -2270
rect 9990 -2390 10002 -2270
rect 9619 -2508 9684 -2406
rect 9619 -4516 9696 -2508
rect 9619 -4618 9684 -4516
rect 9619 -4830 9696 -4618
rect 9814 -4630 10002 -2390
rect 10120 -2406 10197 -2030
rect 10132 -2508 10197 -2406
rect 10120 -4516 10197 -2508
rect 10132 -4618 10197 -4516
rect 9814 -4750 9820 -4630
rect 9990 -4750 10002 -4630
rect 9814 -4770 10002 -4750
rect 10120 -4770 10197 -4618
rect 10229 -1910 10306 -1890
rect 10229 -2030 10230 -1910
rect 10300 -2030 10306 -1910
rect 10229 -2406 10306 -2030
rect 13780 -1910 13857 -1890
rect 13850 -2030 13857 -1910
rect 11340 -2090 11417 -2070
rect 11410 -2210 11417 -2090
rect 10424 -2270 10612 -2250
rect 10424 -2390 10430 -2270
rect 10600 -2390 10612 -2270
rect 10229 -2508 10294 -2406
rect 10229 -4516 10306 -2508
rect 10229 -4618 10294 -4516
rect 10229 -4770 10306 -4618
rect 10424 -4630 10612 -2390
rect 10730 -2406 10807 -2250
rect 10742 -2508 10807 -2406
rect 10730 -4516 10807 -2508
rect 10742 -4618 10807 -4516
rect 10424 -4750 10430 -4630
rect 10600 -4750 10612 -4630
rect 10424 -4770 10612 -4750
rect 10730 -4830 10807 -4618
rect 10839 -2406 10916 -2250
rect 11034 -2270 11222 -2250
rect 11034 -2390 11040 -2270
rect 11210 -2390 11222 -2270
rect 10839 -2508 10904 -2406
rect 10839 -4516 10916 -2508
rect 10839 -4618 10904 -4516
rect 10839 -4830 10916 -4618
rect 11034 -4630 11222 -2390
rect 11340 -2406 11417 -2210
rect 12669 -2090 12746 -2070
rect 12669 -2210 12670 -2090
rect 12740 -2210 12746 -2090
rect 11352 -2508 11417 -2406
rect 11340 -4516 11417 -2508
rect 11352 -4618 11417 -4516
rect 11034 -4750 11040 -4630
rect 11210 -4750 11222 -4630
rect 11034 -4770 11222 -4750
rect 11340 -4770 11417 -4618
rect 11449 -2406 11526 -2250
rect 11644 -2270 11832 -2250
rect 11644 -2390 11650 -2270
rect 11820 -2390 11832 -2270
rect 11449 -2508 11514 -2406
rect 11449 -4516 11526 -2508
rect 11449 -4618 11514 -4516
rect 11449 -4620 11526 -4618
rect 11449 -4630 11530 -4620
rect 11644 -4630 11832 -2390
rect 11950 -2270 12136 -2250
rect 11950 -2390 11960 -2270
rect 12130 -2390 12136 -2270
rect 11950 -2406 12136 -2390
rect 12254 -2270 12442 -2250
rect 12254 -2390 12260 -2270
rect 12430 -2390 12442 -2270
rect 11962 -2508 12124 -2406
rect 11950 -4516 12136 -2508
rect 11962 -4618 12124 -4516
rect 11449 -4770 11600 -4630
rect 11644 -4750 11650 -4630
rect 11820 -4750 11832 -4630
rect 11644 -4770 11832 -4750
rect 11950 -4630 12136 -4618
rect 11950 -4750 11960 -4630
rect 12130 -4750 12136 -4630
rect 11950 -4770 12136 -4750
rect 12254 -4630 12442 -2390
rect 12560 -2406 12637 -2250
rect 12572 -2508 12637 -2406
rect 12560 -4516 12637 -2508
rect 12572 -4618 12637 -4516
rect 12560 -4620 12637 -4618
rect 12254 -4750 12260 -4630
rect 12430 -4750 12442 -4630
rect 12254 -4770 12442 -4750
rect 12490 -4770 12637 -4620
rect 12669 -2406 12746 -2210
rect 12864 -2270 13052 -2250
rect 12864 -2390 12870 -2270
rect 13040 -2390 13052 -2270
rect 12669 -2508 12734 -2406
rect 12669 -4516 12746 -2508
rect 12669 -4618 12734 -4516
rect 12669 -4770 12746 -4618
rect 12864 -4630 13052 -2390
rect 13170 -2406 13247 -2250
rect 13182 -2508 13247 -2406
rect 13170 -4516 13247 -2508
rect 13182 -4618 13247 -4516
rect 12864 -4750 12870 -4630
rect 13040 -4750 13052 -4630
rect 12864 -4770 13052 -4750
rect 11450 -4830 11600 -4770
rect 12490 -4830 12630 -4770
rect 13170 -4830 13247 -4618
rect 13279 -2406 13356 -2250
rect 13474 -2270 13662 -2250
rect 13474 -2390 13480 -2270
rect 13650 -2390 13662 -2270
rect 13279 -2508 13344 -2406
rect 13279 -4516 13356 -2508
rect 13279 -4618 13344 -4516
rect 13279 -4830 13356 -4618
rect 13474 -4630 13662 -2390
rect 13780 -2406 13857 -2030
rect 13792 -2508 13857 -2406
rect 13780 -4516 13857 -2508
rect 13792 -4618 13857 -4516
rect 13474 -4750 13480 -4630
rect 13650 -4750 13662 -4630
rect 13474 -4770 13662 -4750
rect 13780 -4770 13857 -4618
rect 13889 -1910 13966 -1890
rect 13889 -2030 13890 -1910
rect 13960 -2030 13966 -1910
rect 13889 -2406 13966 -2030
rect 15000 -1910 15077 -1890
rect 15070 -2030 15077 -1910
rect 14084 -2270 14272 -2250
rect 14084 -2390 14090 -2270
rect 14260 -2390 14272 -2270
rect 13889 -2508 13954 -2406
rect 13889 -4516 13966 -2508
rect 13889 -4618 13954 -4516
rect 13889 -4770 13966 -4618
rect 14084 -4630 14272 -2390
rect 14390 -2406 14467 -2250
rect 14402 -2508 14467 -2406
rect 14390 -4516 14467 -2508
rect 14402 -4618 14467 -4516
rect 14084 -4750 14090 -4630
rect 14260 -4750 14272 -4630
rect 14084 -4770 14272 -4750
rect 14390 -4830 14467 -4618
rect 14499 -2406 14576 -2250
rect 14694 -2270 14882 -2250
rect 14694 -2390 14700 -2270
rect 14870 -2390 14882 -2270
rect 14499 -2508 14564 -2406
rect 14499 -4516 14576 -2508
rect 14499 -4618 14564 -4516
rect 14499 -4830 14576 -4618
rect 14694 -4630 14882 -2390
rect 15000 -2406 15077 -2030
rect 15012 -2508 15077 -2406
rect 15000 -4516 15077 -2508
rect 15012 -4618 15077 -4516
rect 14694 -4750 14700 -4630
rect 14870 -4750 14882 -4630
rect 14694 -4770 14882 -4750
rect 15000 -4770 15077 -4618
rect 15109 -1910 15186 -1890
rect 15109 -2030 15110 -1910
rect 15180 -2030 15186 -1910
rect 15109 -2406 15186 -2030
rect 15304 -2270 15492 -2250
rect 15304 -2390 15310 -2270
rect 15480 -2390 15492 -2270
rect 15109 -2508 15174 -2406
rect 15109 -4516 15186 -2508
rect 15109 -4618 15174 -4516
rect 15109 -4770 15186 -4618
rect 15304 -4630 15492 -2390
rect 15610 -2406 15687 -2250
rect 15622 -2508 15687 -2406
rect 15610 -4516 15687 -2508
rect 15622 -4618 15687 -4516
rect 15304 -4750 15310 -4630
rect 15480 -4750 15492 -4630
rect 15304 -4770 15492 -4750
rect 15610 -4830 15687 -4618
rect 15719 -2406 15796 -1830
rect 15719 -2508 15784 -2406
rect 15719 -4516 15796 -2508
rect 15719 -4618 15784 -4516
rect 15719 -4830 15796 -4618
rect 15914 -4830 16102 -1830
rect 16220 -1870 16510 -1830
rect 16220 -2406 16380 -1870
rect 16232 -2508 16380 -2406
rect 16220 -4516 16380 -2508
rect 16232 -4618 16380 -4516
rect 16220 -4790 16380 -4618
rect 16430 -4790 16510 -1870
rect 16220 -4830 16510 -4790
rect -1490 -4840 16510 -4830
rect -1490 -4890 -1160 -4840
rect 7410 -4890 7760 -4840
rect 16330 -4890 16510 -4840
rect -1490 -5360 16510 -4890
rect 17240 -6170 17520 -1030
rect 17240 -6390 17250 -6170
rect 17510 -6390 17520 -6170
rect 17240 -6400 17520 -6390
<< via1 >>
rect 2390 8460 2570 8580
rect 2390 6080 2570 6200
rect 2810 8460 2870 8580
rect 3000 8460 3180 8580
rect 2810 6080 2870 6200
rect 3000 6080 3180 6200
rect 3610 8460 3790 8580
rect 3920 8460 3980 8580
rect 3610 6080 3790 6200
rect 3920 6080 3980 6200
rect 4220 8460 4400 8580
rect 2700 5900 2760 6020
rect 4220 6080 4400 6200
rect 4030 5900 4090 6020
rect 8620 8460 8800 8580
rect 8620 6080 8800 6200
rect 8930 5900 8990 6020
rect 9230 8460 9410 8580
rect 9230 6080 9410 6200
rect 9840 8460 10020 8580
rect 9840 6080 10020 6200
rect 9040 5900 9100 6020
rect 10150 5900 10210 6020
rect 10450 8460 10630 8580
rect 10450 6080 10630 6200
rect 11060 8460 11240 8580
rect 11060 6080 11240 6200
rect 10260 5900 10320 6020
rect 11480 8460 11540 8580
rect 11670 8460 11850 8580
rect 11480 6080 11540 6200
rect 11670 6080 11850 6200
rect 12280 8460 12460 8580
rect 12590 8460 12650 8580
rect 12280 6080 12460 6200
rect 12590 6080 12650 6200
rect 12890 8460 13070 8580
rect 11370 5900 11430 6020
rect 12890 6080 13070 6200
rect 13500 8460 13680 8580
rect 13500 6080 13680 6200
rect 12700 5900 12760 6020
rect 13810 5900 13870 6020
rect 14110 8460 14290 8580
rect 13920 5900 13980 6020
rect 14110 6080 14290 6200
rect 14720 8460 14900 8580
rect 14720 6080 14900 6200
rect 15030 5900 15090 6020
rect 15330 8460 15510 8580
rect 15330 6080 15510 6200
rect 15140 5900 15200 6020
rect -230 4380 80 4500
rect -230 10 80 130
rect 1710 4560 1780 4680
rect 1880 10 2090 130
rect 2200 -170 2270 -50
rect 2320 4560 2390 4680
rect 2490 10 2700 130
rect 2810 -170 2880 -50
rect 2930 4740 3000 4860
rect 3100 4380 3310 4500
rect 3420 -350 3490 -230
rect 3540 -170 3610 -50
rect 4030 4560 4100 4680
rect 3710 10 3920 130
rect 4320 4380 4530 4500
rect 4150 -350 4220 -230
rect 4640 4740 4710 4860
rect 4760 4740 4830 4860
rect 4930 4380 5140 4500
rect 5250 -350 5320 -230
rect 5370 4560 5440 4680
rect 5540 10 5750 130
rect 5860 -170 5930 -50
rect 6150 4380 6360 4500
rect 5980 -350 6050 -230
rect 6470 4740 6540 4860
rect 6590 -170 6660 -50
rect 7080 4560 7150 4680
rect 6760 10 6970 130
rect 7370 4380 7580 4500
rect 7200 -350 7270 -230
rect 7690 4740 7760 4860
rect 9880 4930 9960 5050
rect 10190 4930 10270 5050
rect 9880 550 9960 670
rect 10500 4930 10580 5050
rect 10190 550 10270 670
rect 10810 4930 10890 5050
rect 10500 550 10580 670
rect 10010 370 10150 490
rect 11120 4930 11200 5050
rect 10810 550 10890 670
rect 11430 4930 11510 5050
rect 11120 550 11200 670
rect 10630 370 10770 490
rect 11740 4930 11820 5050
rect 11430 550 11510 670
rect 12050 4930 12130 5050
rect 11740 550 11820 670
rect 11250 370 11390 490
rect 12360 4930 12440 5050
rect 12050 550 12130 670
rect 12670 4930 12750 5050
rect 12360 550 12440 670
rect 11870 370 12010 490
rect 12980 4930 13060 5050
rect 12670 550 12750 670
rect 13290 4930 13370 5050
rect 12980 550 13060 670
rect 12490 370 12630 490
rect 13600 4930 13680 5050
rect 13290 550 13370 670
rect 13910 4930 13990 5050
rect 13600 550 13680 670
rect 13110 370 13250 490
rect 14220 4930 14300 5050
rect 13910 550 13990 670
rect 14530 4930 14610 5050
rect 14220 550 14300 670
rect 13730 370 13870 490
rect 14840 4930 14920 5050
rect 14530 550 14610 670
rect 15150 4930 15230 5050
rect 14840 550 14920 670
rect 14350 370 14490 490
rect 15460 4930 15540 5050
rect 15150 550 15230 670
rect 15770 4930 15850 5050
rect 15460 550 15540 670
rect 14970 370 15110 490
rect 15770 550 15850 670
rect 15590 370 15730 490
rect 16700 350 17510 820
rect 9070 -580 9590 -280
rect 11440 -1010 11840 -800
rect 12050 -1010 12450 -800
rect 12670 -1010 13070 -800
rect 13300 -1010 13690 -800
rect 6100 -1550 6640 -1170
rect 7730 -1550 8270 -1170
rect -20 -2210 50 -2090
rect -320 -2390 -150 -2270
rect -320 -4750 -150 -4630
rect 90 -2210 160 -2090
rect 1200 -2210 1270 -2090
rect 290 -2390 460 -2270
rect 290 -4750 460 -4630
rect 900 -2390 1070 -2270
rect 900 -4750 1070 -4630
rect 1310 -2210 1380 -2090
rect 2420 -2210 2490 -2090
rect 1510 -2390 1680 -2270
rect 1510 -4750 1680 -4630
rect 2120 -2390 2290 -2270
rect 3750 -2210 3820 -2090
rect 2120 -4750 2290 -4630
rect 2530 -2390 2600 -2270
rect 2730 -2390 2900 -2270
rect 2530 -4750 2600 -4630
rect 2730 -4750 2900 -4630
rect 3340 -2390 3510 -2270
rect 3640 -2390 3710 -2270
rect 3340 -4750 3510 -4630
rect 3640 -4750 3710 -4630
rect 4860 -2210 4930 -2090
rect 3950 -2390 4120 -2270
rect 3950 -4750 4120 -4630
rect 4560 -2390 4730 -2270
rect 4560 -4750 4730 -4630
rect 4970 -2210 5040 -2090
rect 6080 -2210 6150 -2090
rect 5170 -2390 5340 -2270
rect 5170 -4750 5340 -4630
rect 5780 -2390 5950 -2270
rect 5780 -4750 5950 -4630
rect 6190 -2210 6260 -2090
rect 6390 -2390 6560 -2270
rect 6390 -4750 6560 -4630
rect 8900 -2030 8970 -1910
rect 8600 -2390 8770 -2270
rect 8600 -4750 8770 -4630
rect 9010 -2030 9080 -1910
rect 10120 -2030 10190 -1910
rect 9210 -2390 9380 -2270
rect 9210 -4750 9380 -4630
rect 9820 -2390 9990 -2270
rect 9820 -4750 9990 -4630
rect 10230 -2030 10300 -1910
rect 13780 -2030 13850 -1910
rect 11340 -2210 11410 -2090
rect 10430 -2390 10600 -2270
rect 10430 -4750 10600 -4630
rect 11040 -2390 11210 -2270
rect 12670 -2210 12740 -2090
rect 11040 -4750 11210 -4630
rect 11650 -2390 11820 -2270
rect 11960 -2390 12130 -2270
rect 12260 -2390 12430 -2270
rect 11650 -4750 11820 -4630
rect 11960 -4750 12130 -4630
rect 12260 -4750 12430 -4630
rect 12870 -2390 13040 -2270
rect 12870 -4750 13040 -4630
rect 13480 -2390 13650 -2270
rect 13480 -4750 13650 -4630
rect 13890 -2030 13960 -1910
rect 15000 -2030 15070 -1910
rect 14090 -2390 14260 -2270
rect 14090 -4750 14260 -4630
rect 14700 -2390 14870 -2270
rect 14700 -4750 14870 -4630
rect 15110 -2030 15180 -1910
rect 15310 -2390 15480 -2270
rect 15310 -4750 15480 -4630
rect 17250 -6390 17510 -6170
<< metal2 >>
rect 1570 8580 5230 8590
rect 1570 8460 2390 8580
rect 2570 8460 2810 8580
rect 2870 8460 3000 8580
rect 3180 8460 3610 8580
rect 3790 8460 3920 8580
rect 3980 8460 4220 8580
rect 4400 8460 5230 8580
rect 1570 8450 5230 8460
rect 7810 8580 16330 8590
rect 7810 8460 8620 8580
rect 8800 8460 9230 8580
rect 9410 8460 9840 8580
rect 10020 8460 10450 8580
rect 10630 8460 11060 8580
rect 11240 8460 11480 8580
rect 11540 8460 11670 8580
rect 11850 8460 12280 8580
rect 12460 8460 12590 8580
rect 12650 8460 12890 8580
rect 13070 8460 13500 8580
rect 13680 8460 14110 8580
rect 14290 8460 14720 8580
rect 14900 8460 15330 8580
rect 15510 8460 16330 8580
rect 7810 8450 16330 8460
rect 1570 6200 7660 6210
rect 1570 6080 2390 6200
rect 2570 6080 2810 6200
rect 2870 6080 3000 6200
rect 3180 6080 3610 6200
rect 3790 6080 3920 6200
rect 3980 6080 4220 6200
rect 4400 6080 7660 6200
rect 1570 6070 7660 6080
rect -860 6020 5230 6030
rect -860 5900 2700 6020
rect 2760 5900 4030 6020
rect 4090 5900 5230 6020
rect -860 5890 5230 5900
rect -860 -2260 -380 5890
rect 7270 4870 7660 6070
rect 7810 6200 16330 6210
rect 7810 6080 8620 6200
rect 8800 6080 9230 6200
rect 9410 6080 9840 6200
rect 10020 6080 10450 6200
rect 10630 6080 11060 6200
rect 11240 6080 11480 6200
rect 11540 6080 11670 6200
rect 11850 6080 12280 6200
rect 12460 6080 12590 6200
rect 12650 6080 12890 6200
rect 13070 6080 13500 6200
rect 13680 6080 14110 6200
rect 14290 6080 14720 6200
rect 14900 6080 15330 6200
rect 15510 6080 16330 6200
rect 7810 6070 16330 6080
rect 1270 4860 7770 4870
rect 1270 4740 2930 4860
rect 3000 4740 4640 4860
rect 4710 4740 4760 4860
rect 4830 4740 6470 4860
rect 6540 4740 7690 4860
rect 7760 4740 7770 4860
rect 1270 4730 7770 4740
rect 7810 4690 8200 6070
rect 8910 6020 16410 6030
rect 8910 5900 8930 6020
rect 8990 5900 9040 6020
rect 9100 5900 10150 6020
rect 10210 5900 10260 6020
rect 10320 5900 11370 6020
rect 11430 5900 12700 6020
rect 12760 5900 13810 6020
rect 13870 5900 13920 6020
rect 13980 5900 15030 6020
rect 15090 5900 15140 6020
rect 15200 5900 16410 6020
rect 8910 5890 16410 5900
rect 1270 4680 8200 4690
rect 1270 4560 1710 4680
rect 1780 4560 2320 4680
rect 2390 4560 4030 4680
rect 4100 4560 5370 4680
rect 5440 4560 7080 4680
rect 7150 4560 8200 4680
rect 1270 4550 8200 4560
rect 9060 5060 9600 5890
rect 16010 5060 16410 5890
rect 9060 5050 16410 5060
rect 9060 4930 9880 5050
rect 9960 4930 10190 5050
rect 10270 4930 10500 5050
rect 10580 4930 10810 5050
rect 10890 4930 11120 5050
rect 11200 4930 11430 5050
rect 11510 4930 11740 5050
rect 11820 4930 12050 5050
rect 12130 4930 12360 5050
rect 12440 4930 12670 5050
rect 12750 4930 12980 5050
rect 13060 4930 13290 5050
rect 13370 4930 13600 5050
rect 13680 4930 13910 5050
rect 13990 4930 14220 5050
rect 14300 4930 14530 5050
rect 14610 4930 14840 5050
rect 14920 4930 15150 5050
rect 15230 4930 15460 5050
rect 15540 4930 15770 5050
rect 15850 4930 16410 5050
rect 9060 4920 16410 4930
rect -240 4500 8430 4510
rect -240 4380 -230 4500
rect 80 4380 3100 4500
rect 3310 4380 4320 4500
rect 4530 4380 4930 4500
rect 5140 4380 6150 4500
rect 6360 4380 7370 4500
rect 7580 4380 8430 4500
rect -240 4370 8430 4380
rect 9060 680 9600 4920
rect 16010 680 16410 4920
rect 9060 670 16410 680
rect 9060 550 9880 670
rect 9960 550 10190 670
rect 10270 550 10500 670
rect 10580 550 10810 670
rect 10890 550 11120 670
rect 11200 550 11430 670
rect 11510 550 11740 670
rect 11820 550 12050 670
rect 12130 550 12360 670
rect 12440 550 12670 670
rect 12750 550 12980 670
rect 13060 550 13290 670
rect 13370 550 13600 670
rect 13680 550 13910 670
rect 13990 550 14220 670
rect 14300 550 14530 670
rect 14610 550 14840 670
rect 14920 550 15150 670
rect 15230 550 15460 670
rect 15540 550 15770 670
rect 15850 550 16410 670
rect 9060 540 16410 550
rect 16690 1340 17520 1350
rect 16690 840 16700 1340
rect 17510 840 17520 1340
rect 16690 820 17520 840
rect -240 130 8430 140
rect -240 10 -230 130
rect 80 10 1880 130
rect 2090 10 2490 130
rect 2700 10 3710 130
rect 3920 10 5540 130
rect 5750 10 6760 130
rect 6970 10 8430 130
rect -240 0 8430 10
rect 1270 -50 8430 -40
rect 1270 -170 2200 -50
rect 2270 -170 2810 -50
rect 2880 -170 3540 -50
rect 3610 -170 5860 -50
rect 5930 -170 6590 -50
rect 6660 -170 8430 -50
rect 1270 -230 8430 -170
rect 1270 -350 3420 -230
rect 3490 -350 4150 -230
rect 4220 -350 5250 -230
rect 5320 -350 5980 -230
rect 6050 -350 7200 -230
rect 7270 -350 8430 -230
rect 1270 -360 8430 -350
rect 9060 -280 9600 540
rect 9770 490 16090 500
rect 9770 370 10010 490
rect 10150 370 10630 490
rect 10770 370 11250 490
rect 11390 370 11870 490
rect 12010 370 12490 490
rect 12630 370 13110 490
rect 13250 370 13730 490
rect 13870 370 14350 490
rect 14490 370 14970 490
rect 15110 370 15590 490
rect 15730 370 16090 490
rect 9770 200 16090 370
rect 16690 350 16700 820
rect 17510 350 17520 820
rect 16690 340 17520 350
rect 6090 -1170 6650 -360
rect 9060 -580 9070 -280
rect 9590 -580 9600 -280
rect 9060 -590 9600 -580
rect 6090 -1550 6100 -1170
rect 6640 -1550 6650 -1170
rect 6090 -1560 6650 -1550
rect 6950 -1060 9600 -590
rect 11420 -800 11840 200
rect 11420 -1010 11440 -800
rect 6950 -2080 7520 -1060
rect -30 -2090 7520 -2080
rect -30 -2210 -20 -2090
rect 50 -2210 90 -2090
rect 160 -2210 1200 -2090
rect 1270 -2210 1310 -2090
rect 1380 -2210 2420 -2090
rect 2490 -2210 3750 -2090
rect 3820 -2210 4860 -2090
rect 4930 -2210 4970 -2090
rect 5040 -2210 6080 -2090
rect 6150 -2210 6190 -2090
rect 6260 -2210 7520 -2090
rect -30 -2220 7520 -2210
rect 7720 -1170 8300 -1160
rect 7720 -1550 7730 -1170
rect 8270 -1550 8300 -1170
rect 7720 -2080 8300 -1550
rect 11420 -1690 11840 -1010
rect 12040 -800 12460 200
rect 12040 -1010 12050 -800
rect 12450 -1010 12460 -800
rect 12040 -1690 12460 -1010
rect 12660 -800 13080 200
rect 12660 -1010 12670 -800
rect 13070 -1010 13080 -800
rect 12660 -1690 13080 -1010
rect 13280 -800 13700 200
rect 13280 -1010 13300 -800
rect 13690 -1010 13700 -800
rect 13280 -1630 13700 -1010
rect 13280 -1690 17170 -1630
rect 11420 -1900 17170 -1690
rect 8890 -1910 17170 -1900
rect 8890 -2030 8900 -1910
rect 8970 -2030 9010 -1910
rect 9080 -2030 10120 -1910
rect 10190 -2030 10230 -1910
rect 10300 -2030 13780 -1910
rect 13850 -2030 13890 -1910
rect 13960 -2030 15000 -1910
rect 15070 -2030 15110 -1910
rect 15180 -2030 17170 -1910
rect 8890 -2040 17170 -2030
rect 7720 -2090 16440 -2080
rect 7720 -2210 11340 -2090
rect 11410 -2210 12670 -2090
rect 12740 -2210 16440 -2090
rect 7720 -2220 16440 -2210
rect -860 -2270 7520 -2260
rect -860 -2390 -320 -2270
rect -150 -2390 290 -2270
rect 460 -2390 900 -2270
rect 1070 -2390 1510 -2270
rect 1680 -2390 2120 -2270
rect 2290 -2390 2530 -2270
rect 2600 -2390 2730 -2270
rect 2900 -2390 3340 -2270
rect 3510 -2390 3640 -2270
rect 3710 -2390 3950 -2270
rect 4120 -2390 4560 -2270
rect 4730 -2390 5170 -2270
rect 5340 -2390 5780 -2270
rect 5950 -2390 6390 -2270
rect 6560 -2390 7520 -2270
rect -860 -2400 7520 -2390
rect 7720 -2270 16440 -2260
rect 7720 -2390 8600 -2270
rect 8770 -2390 9210 -2270
rect 9380 -2390 9820 -2270
rect 9990 -2390 10430 -2270
rect 10600 -2390 11040 -2270
rect 11210 -2390 11650 -2270
rect 11820 -2390 11960 -2270
rect 12130 -2390 12260 -2270
rect 12430 -2390 12870 -2270
rect 13040 -2390 13480 -2270
rect 13650 -2390 14090 -2270
rect 14260 -2390 14700 -2270
rect 14870 -2390 15310 -2270
rect 15480 -2390 16440 -2270
rect 7720 -2400 16440 -2390
rect 16570 -2740 17170 -2040
rect -1200 -4630 7520 -4620
rect -1200 -4750 -320 -4630
rect -150 -4750 290 -4630
rect 460 -4750 900 -4630
rect 1070 -4750 1510 -4630
rect 1680 -4750 2120 -4630
rect 2290 -4750 2530 -4630
rect 2600 -4750 2730 -4630
rect 2900 -4750 3340 -4630
rect 3510 -4750 3640 -4630
rect 3710 -4750 3950 -4630
rect 4120 -4750 4560 -4630
rect 4730 -4750 5170 -4630
rect 5340 -4750 5780 -4630
rect 5950 -4750 6390 -4630
rect 6560 -4750 7520 -4630
rect -1200 -4760 7520 -4750
rect 7720 -4630 15510 -4620
rect 7720 -4750 8600 -4630
rect 8770 -4750 9210 -4630
rect 9380 -4750 9820 -4630
rect 9990 -4750 10430 -4630
rect 10600 -4750 11040 -4630
rect 11210 -4750 11650 -4630
rect 11820 -4750 11960 -4630
rect 12130 -4750 12260 -4630
rect 12430 -4750 12870 -4630
rect 13040 -4750 13480 -4630
rect 13650 -4750 14090 -4630
rect 14260 -4750 14700 -4630
rect 14870 -4750 15310 -4630
rect 15480 -4750 15510 -4630
rect 7720 -4760 15510 -4750
rect 11950 -4830 12140 -4760
rect 7720 -4840 12140 -4830
rect -1490 -5360 12140 -4840
rect -1490 -5910 -780 -5360
rect 17240 -6170 17520 -6160
rect 17240 -6390 17250 -6170
rect 17510 -6390 17520 -6170
rect 17240 -6410 17520 -6390
rect 17240 -6800 17250 -6410
rect 17510 -6800 17520 -6410
rect 17240 -6810 17520 -6800
<< via2 >>
rect 16700 840 17510 1340
rect 17250 -6800 17510 -6410
<< metal3 >>
rect 16690 1800 17520 1810
rect 16690 1360 16700 1800
rect 17510 1360 17520 1800
rect 16690 1340 17520 1360
rect 16690 840 16700 1340
rect 17510 840 17520 1340
rect 16690 830 17520 840
rect 17240 -6410 17520 -6400
rect 17240 -6800 17250 -6410
rect 17510 -6800 17520 -6410
rect 17240 -6820 17520 -6800
rect 17240 -7200 17250 -6820
rect 17510 -7200 17520 -6820
rect 17240 -7210 17520 -7200
<< via3 >>
rect 16700 1360 17510 1800
rect 17250 -7200 17510 -6820
<< metal4 >>
rect -758 8771 17521 9150
rect 1294 -8259 1504 8481
rect 3494 -8169 3704 8771
rect 12074 8770 17521 8771
rect 5694 -8259 5904 8481
rect 9884 -8259 10094 8481
rect 12074 -8169 12284 8770
rect 14264 -8259 14474 8481
rect 16690 1800 17520 8770
rect 16690 1360 16700 1800
rect 17510 1360 17520 1800
rect 16690 1350 17520 1360
rect 1294 -8260 14474 -8259
rect 17240 -6820 17520 -6810
rect 17240 -7200 17250 -6820
rect 17510 -7200 17520 -6820
rect 17240 -8260 17520 -7200
rect 1294 -8479 17520 -8260
rect 17240 -8480 17520 -8479
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_0
timestamp 1650738325
transform 1 0 1454 0 1 6521
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_1
timestamp 1650738325
transform -1 0 5743 0 -1 6521
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_2
timestamp 1650738325
transform -1 0 14323 0 -1 6521
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_3
timestamp 1650738325
transform 1 0 10034 0 1 6521
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_4
timestamp 1650738325
transform -1 0 14323 0 -1 2321
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_5
timestamp 1650738325
transform 1 0 10034 0 1 2321
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_6
timestamp 1650738325
transform 1 0 1454 0 1 2321
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_7
timestamp 1650738325
transform -1 0 5743 0 -1 2321
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_8
timestamp 1650738325
transform -1 0 14323 0 -1 -1879
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_9
timestamp 1650738325
transform 1 0 10034 0 1 -1879
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_10
timestamp 1650738325
transform 1 0 1454 0 1 -1879
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_11
timestamp 1650738325
transform -1 0 5743 0 -1 -1879
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_12
timestamp 1650738325
transform -1 0 14323 0 -1 -6079
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_13
timestamp 1650738325
transform 1 0 10034 0 1 -6079
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_14
timestamp 1650738325
transform 1 0 1454 0 1 -6079
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_15
timestamp 1650738325
transform -1 0 5743 0 -1 -6079
box -2150 -2100 2149 2100
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_0
timestamp 1650752648
transform 1 0 -842 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_1
timestamp 1650752648
transform 1 0 -232 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_2
timestamp 1650752648
transform 1 0 378 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_3
timestamp 1650752648
transform 1 0 988 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_4
timestamp 1650752648
transform 1 0 1598 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_5
timestamp 1650752648
transform 1 0 2208 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_6
timestamp 1650752648
transform 1 0 2818 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_7
timestamp 1650752648
transform 1 0 3428 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_8
timestamp 1650752648
transform 1 0 4038 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_9
timestamp 1650752648
transform 1 0 4648 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_10
timestamp 1650752648
transform 1 0 5258 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_11
timestamp 1650752648
transform 1 0 5868 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_12
timestamp 1650752648
transform 1 0 6478 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_13
timestamp 1650752648
transform 1 0 7088 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_14
timestamp 1650752648
transform 1 0 14788 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_15
timestamp 1650752648
transform 1 0 15398 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_16
timestamp 1650752648
transform 1 0 16008 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_17
timestamp 1650752648
transform 1 0 12958 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_18
timestamp 1650752648
transform 1 0 13568 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_19
timestamp 1650752648
transform 1 0 14178 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_20
timestamp 1650752648
transform 1 0 11738 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_21
timestamp 1650752648
transform 1 0 12348 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_22
timestamp 1650752648
transform 1 0 9908 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_23
timestamp 1650752648
transform 1 0 10518 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_24
timestamp 1650752648
transform 1 0 11128 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_25
timestamp 1650752648
transform 1 0 8078 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_26
timestamp 1650752648
transform 1 0 8688 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_64LW2M  sky130_fd_pr__nfet_g5v0d10v5_64LW2M_27
timestamp 1650752648
transform 1 0 9298 0 1 -3512
box -258 -1088 258 1088
use sky130_fd_pr__nfet_g5v0d10v5_NKLCM2  sky130_fd_pr__nfet_g5v0d10v5_NKLCM2_0
timestamp 1650752648
transform 1 0 1988 0 1 2258
box -258 -2088 258 2088
use sky130_fd_pr__nfet_g5v0d10v5_NKLCM2  sky130_fd_pr__nfet_g5v0d10v5_NKLCM2_1
timestamp 1650752648
transform 1 0 2598 0 1 2258
box -258 -2088 258 2088
use sky130_fd_pr__nfet_g5v0d10v5_NKLCM2  sky130_fd_pr__nfet_g5v0d10v5_NKLCM2_2
timestamp 1650752648
transform 1 0 3208 0 1 2258
box -258 -2088 258 2088
use sky130_fd_pr__nfet_g5v0d10v5_NKLCM2  sky130_fd_pr__nfet_g5v0d10v5_NKLCM2_3
timestamp 1650752648
transform 1 0 3818 0 1 2258
box -258 -2088 258 2088
use sky130_fd_pr__nfet_g5v0d10v5_NKLCM2  sky130_fd_pr__nfet_g5v0d10v5_NKLCM2_4
timestamp 1650752648
transform 1 0 4428 0 1 2258
box -258 -2088 258 2088
use sky130_fd_pr__nfet_g5v0d10v5_NKLCM2  sky130_fd_pr__nfet_g5v0d10v5_NKLCM2_5
timestamp 1650752648
transform 1 0 5038 0 1 2258
box -258 -2088 258 2088
use sky130_fd_pr__nfet_g5v0d10v5_NKLCM2  sky130_fd_pr__nfet_g5v0d10v5_NKLCM2_6
timestamp 1650752648
transform 1 0 5648 0 1 2258
box -258 -2088 258 2088
use sky130_fd_pr__nfet_g5v0d10v5_NKLCM2  sky130_fd_pr__nfet_g5v0d10v5_NKLCM2_7
timestamp 1650752648
transform 1 0 6258 0 1 2258
box -258 -2088 258 2088
use sky130_fd_pr__nfet_g5v0d10v5_NKLCM2  sky130_fd_pr__nfet_g5v0d10v5_NKLCM2_8
timestamp 1650752648
transform 1 0 6868 0 1 2258
box -258 -2088 258 2088
use sky130_fd_pr__nfet_g5v0d10v5_NKLCM2  sky130_fd_pr__nfet_g5v0d10v5_NKLCM2_9
timestamp 1650752648
transform 1 0 7478 0 1 2258
box -258 -2088 258 2088
use sky130_fd_pr__nfet_g5v0d10v5_NKLCM2  sky130_fd_pr__nfet_g5v0d10v5_NKLCM2_10
timestamp 1650752648
transform 1 0 8088 0 1 2258
box -258 -2088 258 2088
use sky130_fd_pr__nfet_g5v0d10v5_NKLCM2  sky130_fd_pr__nfet_g5v0d10v5_NKLCM2_11
timestamp 1650752648
transform 1 0 1378 0 1 2258
box -258 -2088 258 2088
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_4
timestamp 1649000094
transform 1 0 1874 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_5
timestamp 1649000094
transform 1 0 2484 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_6
timestamp 1649000094
transform 1 0 3094 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_7
timestamp 1649000094
transform 1 0 3704 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_8
timestamp 1649000094
transform 1 0 4314 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_9
timestamp 1649000094
transform 1 0 4924 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_14
timestamp 1649000094
transform 1 0 15424 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_15
timestamp 1649000094
transform 1 0 16034 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_16
timestamp 1649000094
transform 1 0 13594 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_17
timestamp 1649000094
transform 1 0 14204 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_18
timestamp 1649000094
transform 1 0 14814 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_19
timestamp 1649000094
transform 1 0 12374 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_20
timestamp 1649000094
transform 1 0 12984 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_21
timestamp 1649000094
transform 1 0 10544 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_22
timestamp 1649000094
transform 1 0 11154 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_23
timestamp 1649000094
transform 1 0 11764 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_24
timestamp 1649000094
transform 1 0 9324 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_25
timestamp 1649000094
transform 1 0 9934 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_26
timestamp 1649000094
transform 1 0 8104 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_PCRJQC  sky130_fd_pr__pfet_g5v0d10v5_PCRJQC_27
timestamp 1649000094
transform 1 0 8714 0 1 7330
box -324 -1100 324 1100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_0
timestamp 1650751748
transform 1 0 9924 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_1
timestamp 1650751748
transform 1 0 10234 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_2
timestamp 1650751748
transform 1 0 10544 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_3
timestamp 1650751748
transform 1 0 10854 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_4
timestamp 1650751748
transform 1 0 11164 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_5
timestamp 1650751748
transform 1 0 11474 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_6
timestamp 1650751748
transform 1 0 11784 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_7
timestamp 1650751748
transform 1 0 12094 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_8
timestamp 1650751748
transform 1 0 12404 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_9
timestamp 1650751748
transform 1 0 12714 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_10
timestamp 1650751748
transform 1 0 13024 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_11
timestamp 1650751748
transform 1 0 13334 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_12
timestamp 1650751748
transform 1 0 13644 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_13
timestamp 1650751748
transform 1 0 13954 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_14
timestamp 1650751748
transform 1 0 14264 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_15
timestamp 1650751748
transform 1 0 14574 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_16
timestamp 1650751748
transform 1 0 14884 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_17
timestamp 1650751748
transform 1 0 15194 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_18
timestamp 1650751748
transform 1 0 15504 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD  sky130_fd_pr__pfet_g5v0d10v5_Y6SSWD_19
timestamp 1650751748
transform 1 0 15814 0 1 2800
box -174 -2100 174 2100
use sky130_fd_pr__res_xhigh_po_1p41_YMGX8A  sky130_fd_pr__res_xhigh_po_1p41_YMGX8A_0
timestamp 1725111857
transform 0 1 15162 -1 0 -1323
box -307 -782 307 782
<< labels >>
flabel metal1 -1490 0 -990 700 0 FreeSans 1600 0 0 0 INN
port 4 nsew
flabel metal1 -1490 3810 -990 4510 0 FreeSans 1600 0 0 0 INP
port 5 nsew
flabel metal1 -1490 5450 -1090 9150 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal1 -1490 -1770 -990 -370 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal2 -1490 -5910 -780 -5050 0 FreeSans 1600 0 0 0 IB
port 3 nsew
flabel metal2 16570 -2740 17170 -1630 0 FreeSans 1600 0 0 0 VOUT
port 2 nsew
<< end >>
