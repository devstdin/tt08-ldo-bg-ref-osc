magic
tech sky130A
magscale 1 2
timestamp 1725192368
<< nwell >>
rect -3331 12250 -148 12255
rect -3331 11539 6450 12250
rect -3332 9220 6450 11539
rect -3332 9175 2600 9220
rect -3332 9174 -109 9175
rect -3332 6823 -542 9174
<< mvnsubdiff >>
rect 710 12090 5810 12130
rect 710 11990 750 12090
rect 5770 11990 5810 12090
rect 710 11950 5810 11990
rect 6190 11730 6360 11770
rect 100 11590 510 11620
rect -792 11427 -642 11467
rect -792 6930 -752 11427
rect -672 6930 -642 11427
rect 100 9680 130 11590
rect 480 9680 510 11590
rect 6190 10390 6230 11730
rect 6320 10390 6360 11730
rect 6190 10350 6360 10390
rect 100 9650 510 9680
rect 860 9410 5200 9440
rect 860 9320 900 9410
rect 5160 9320 5200 9410
rect 860 9290 5200 9320
rect -792 6907 -642 6930
<< mvnsubdiffcont >>
rect 750 11990 5770 12090
rect -752 6930 -672 11427
rect 130 9680 480 11590
rect 6230 10390 6320 11730
rect 900 9320 5160 9410
<< locali >>
rect 730 12090 5790 12110
rect 730 11990 750 12090
rect 5770 11990 5790 12090
rect 730 11970 5790 11990
rect 6210 11730 6340 11750
rect 110 11590 500 11610
rect -772 11427 -662 11447
rect -772 6930 -752 11427
rect -672 6930 -662 11427
rect 110 9680 130 11590
rect 480 9680 500 11590
rect 6210 10390 6230 11730
rect 6320 10390 6340 11730
rect 6210 10370 6340 10390
rect 110 9660 500 9680
rect 880 9410 5180 9430
rect 880 9320 900 9410
rect 5160 9320 5180 9410
rect 880 9300 5180 9320
rect -772 6914 -662 6930
rect 740 3600 1860 3730
rect 740 2760 880 3600
rect 1720 2760 1860 3600
rect 740 2650 1860 2760
rect 1090 2620 1860 2650
rect 2030 3600 3150 3730
rect 2030 2760 2170 3600
rect 3010 2760 3150 3600
rect 2030 2650 3150 2760
rect 3320 3600 4430 3730
rect 3320 2760 3460 3600
rect 4300 2760 4430 3600
rect 3320 2650 4430 2760
rect 2030 2620 2250 2650
rect 1090 2420 1860 2440
rect 740 2310 1860 2420
rect 740 1470 880 2310
rect 1720 1470 1860 2310
rect 740 1360 1860 1470
rect 2030 2420 2250 2440
rect 3420 2620 4080 2650
rect 3420 2420 4080 2440
rect 2030 2310 3120 2420
rect 2030 1470 2170 2310
rect 3010 1470 3120 2310
rect 2030 1360 3120 1470
rect 3350 2310 4430 2420
rect 3350 1470 3460 2310
rect 4300 1470 4430 2310
rect 3350 1360 4430 1470
rect 1090 1330 1770 1360
rect 1090 1130 1770 1160
rect 3420 1330 4080 1360
rect 3420 1130 4080 1160
rect 740 1020 1860 1130
rect 740 180 880 1020
rect 1720 420 1860 1020
rect 2030 1020 3150 1130
rect 2030 420 2170 1020
rect 1720 180 1830 420
rect 740 40 1830 180
rect 2060 180 2170 420
rect 3010 420 3150 1020
rect 3320 1020 4430 1130
rect 3320 420 3460 1020
rect 3010 180 3120 420
rect 2060 40 3120 180
rect 3350 180 3460 420
rect 4300 180 4430 1020
rect 3350 40 4430 180
rect 4960 1060 6090 1210
rect 4960 220 5100 1060
rect 5950 220 6090 1060
rect 4960 80 6090 220
<< viali >>
rect 750 11990 5770 12090
rect -752 6930 -672 11427
rect 130 9680 480 11590
rect 6230 10390 6320 11730
rect 900 9320 5160 9410
rect -52 8103 -18 8453
rect 2406 8103 2440 8453
rect -52 7595 -18 7945
rect 4890 7440 4924 7790
rect -52 7087 -18 7437
rect 2406 7087 2440 7437
rect -2695 6720 -2489 6754
rect -2331 6720 -2125 6754
rect -1967 6720 -1761 6754
rect -1603 6720 -1397 6754
rect -1239 6720 -1033 6754
rect -875 6720 -669 6754
rect -52 6579 -18 6929
rect 2406 6579 2440 6929
rect 4890 6910 4924 7260
rect 3024 6694 3374 6728
rect 3532 6694 3882 6728
rect 4040 6694 4390 6728
rect -52 6071 -18 6421
rect 2406 6071 2440 6421
rect 4890 6380 4924 6730
rect -52 5563 -18 5913
rect 2406 5563 2440 5913
rect 4890 5850 4924 6200
rect -52 5055 -18 5405
rect 4890 5320 4924 5670
rect -52 4547 -18 4897
rect 2406 4547 2440 4897
rect 4890 4790 4924 5140
rect 3024 4236 3374 4270
rect 4040 4236 4390 4270
rect 4890 4260 4924 4610
rect 670 3750 1760 3800
rect 2130 3750 3050 3800
rect 3420 3750 4500 3800
rect 670 2650 720 3750
rect 670 2420 1090 2650
rect 4450 2650 4500 3750
rect 4890 3730 4924 4080
rect 4890 3200 4924 3550
rect 4890 2670 4924 3020
rect 670 1360 720 2420
rect 2250 2420 3420 2650
rect 4080 2420 4500 2650
rect 3120 1360 3350 2420
rect 4450 1360 4500 2420
rect 4890 2140 4924 2490
rect 4890 1610 4924 1960
rect 670 1130 1090 1360
rect 1770 1130 3420 1360
rect 4080 1130 4500 1360
rect 670 20 720 1130
rect 1830 20 2060 420
rect 3120 20 3350 420
rect 4450 20 4500 1130
rect 670 -20 4500 20
rect -3059 -138 -2853 -104
rect -2695 -138 -2489 -104
rect -2331 -138 -2125 -104
rect -1967 -138 -1761 -104
rect -1603 -138 -1397 -104
rect -1239 -138 -1033 -104
rect -875 -138 -669 -104
<< metal1 >>
rect -3701 12090 7950 12640
rect -3701 11990 750 12090
rect 5770 11990 7950 12090
rect -3701 11790 7950 11990
rect -3701 11770 1100 11790
rect -3701 11740 550 11770
rect -3701 11602 -3087 11740
rect -907 11602 550 11740
rect -3701 11590 550 11602
rect -3701 11491 130 11590
rect -3701 11427 -582 11491
rect -2972 11387 -2882 11397
rect -2972 11277 -2962 11387
rect -2892 11277 -2882 11387
rect -2972 11267 -2882 11277
rect -3062 11187 -2962 11227
rect -3701 11065 -3072 11137
rect -3701 7061 -3405 11065
rect -3356 7137 -3072 11065
rect -3356 7061 -3142 7137
rect -3032 7097 -2992 11187
rect -2932 11157 -2882 11267
rect -2952 7147 -2882 11157
rect -2852 11267 -2782 11427
rect -2722 11387 -2622 11397
rect -2722 11277 -2712 11387
rect -2632 11277 -2622 11387
rect -2852 11157 -2802 11267
rect -2722 11227 -2622 11277
rect -2462 11267 -2392 11427
rect -2332 11387 -2232 11397
rect -2332 11277 -2322 11387
rect -2242 11277 -2232 11387
rect -2772 11187 -2572 11227
rect -2852 7147 -2782 11157
rect -2722 7097 -2622 11187
rect -2462 11157 -2412 11267
rect -2332 11227 -2232 11277
rect -2072 11267 -2002 11427
rect -1952 11387 -1852 11397
rect -1952 11277 -1942 11387
rect -1862 11277 -1852 11387
rect -2382 11187 -2192 11227
rect -2562 7137 -2492 11137
rect -2462 7147 -2392 11157
rect -3701 -95 -3142 7061
rect -3062 7057 -2962 7097
rect -2762 7057 -2572 7097
rect -3032 7027 -2992 7057
rect -2542 7027 -2492 7137
rect -2332 7097 -2232 11187
rect -2072 11157 -2022 11267
rect -1952 11227 -1852 11277
rect -1692 11267 -1622 11427
rect -1562 11387 -1462 11397
rect -1562 11277 -1552 11387
rect -1472 11277 -1462 11387
rect -1992 11187 -1802 11227
rect -2182 7137 -2112 11137
rect -2072 7147 -2002 11157
rect -2382 7057 -2192 7097
rect -2152 7027 -2112 7137
rect -1952 7097 -1852 11187
rect -1692 11157 -1642 11267
rect -1562 11227 -1462 11277
rect -1302 11267 -1232 11427
rect -1172 11387 -1072 11397
rect -1172 11277 -1162 11387
rect -1082 11277 -1072 11387
rect -1602 11187 -1412 11227
rect -1792 7137 -1722 11137
rect -1692 7147 -1622 11157
rect -1992 7057 -1802 7097
rect -1772 7027 -1722 7137
rect -1562 7097 -1462 11187
rect -1302 11157 -1252 11267
rect -1172 11227 -1072 11277
rect -1212 11187 -1022 11227
rect -1402 7137 -1332 11137
rect -1302 7147 -1232 11157
rect -1602 7057 -1412 7097
rect -1382 7027 -1332 7137
rect -1172 7097 -1072 11187
rect -1012 7137 -932 11157
rect -1212 7057 -1022 7097
rect -992 7027 -932 7137
rect -3032 6937 -932 7027
rect -3032 6197 -2897 6937
rect -812 6930 -752 11427
rect -672 6930 -582 11427
rect 70 9680 130 11491
rect 480 9680 550 11590
rect 650 11400 1100 11770
rect 1160 11720 1250 11730
rect 1160 11410 1170 11720
rect 1240 11410 1250 11720
rect 650 11370 860 11400
rect 650 11290 910 11370
rect 650 10380 710 11290
rect 770 10270 860 11290
rect 950 11260 1080 11400
rect 1160 11370 1250 11410
rect 1550 11720 1640 11730
rect 1550 11410 1560 11720
rect 1630 11410 1640 11720
rect 1550 11370 1640 11410
rect 1710 11400 1870 11790
rect 1940 11720 2030 11730
rect 1940 11410 1950 11720
rect 2020 11410 2030 11720
rect 1110 11290 1300 11370
rect 1500 11290 1690 11370
rect 930 10370 1100 11260
rect 1160 10270 1250 11290
rect 1320 10300 1380 11190
rect 720 10190 910 10270
rect 1110 10190 1300 10270
rect 1330 10160 1380 10300
rect 70 9470 550 9680
rect 1240 9710 1380 10160
rect 1240 9560 1250 9710
rect 1370 9560 1380 9710
rect 1240 9550 1380 9560
rect 1420 10300 1480 11190
rect 1420 10160 1470 10300
rect 1550 10270 1640 11290
rect 1730 11260 1850 11400
rect 1940 11370 2030 11410
rect 2320 11720 2410 11730
rect 2320 11410 2330 11720
rect 2400 11410 2410 11720
rect 2320 11370 2410 11410
rect 2480 11400 2650 11790
rect 2710 11720 2800 11730
rect 2710 11410 2720 11720
rect 2790 11410 2800 11720
rect 1880 11290 2070 11370
rect 2280 11290 2470 11370
rect 1710 10370 1870 11260
rect 1940 10270 2030 11290
rect 2090 10300 2150 11190
rect 1500 10190 1690 10270
rect 1890 10190 2080 10270
rect 2110 10160 2150 10300
rect 1420 9930 1560 10160
rect 1420 9780 1430 9930
rect 1550 9780 1560 9930
rect 1420 9550 1560 9780
rect 2010 10150 2150 10160
rect 2010 10000 2020 10150
rect 2140 10000 2150 10150
rect 2010 9550 2150 10000
rect 2200 10300 2260 11190
rect 2200 10160 2240 10300
rect 2320 10270 2410 11290
rect 2500 11260 2630 11400
rect 2710 11370 2800 11410
rect 3100 11720 3190 11730
rect 3100 11410 3110 11720
rect 3180 11410 3190 11720
rect 3100 11370 3190 11410
rect 3260 11400 3420 11790
rect 3490 11720 3580 11730
rect 3490 11410 3500 11720
rect 3570 11410 3580 11720
rect 2670 11290 2860 11370
rect 3050 11290 3240 11370
rect 2480 10370 2650 11260
rect 2710 10270 2800 11290
rect 2870 10300 2930 11190
rect 2270 10190 2460 10270
rect 2660 10190 2850 10270
rect 2890 10160 2930 10300
rect 2200 9710 2340 10160
rect 2200 9560 2210 9710
rect 2330 9560 2340 9710
rect 2200 9550 2340 9560
rect 2790 9930 2930 10160
rect 2790 9780 2800 9930
rect 2920 9780 2930 9930
rect 2790 9550 2930 9780
rect 2970 10300 3030 11190
rect 2970 10160 3020 10300
rect 3100 10270 3190 11290
rect 3280 11260 3400 11400
rect 3490 11370 3580 11410
rect 3880 11720 3970 11730
rect 3880 11410 3890 11720
rect 3960 11410 3970 11720
rect 3880 11370 3970 11410
rect 4030 11400 4200 11790
rect 4260 11720 4350 11730
rect 4260 11410 4270 11720
rect 4340 11410 4350 11720
rect 3440 11290 3630 11370
rect 3830 11290 4020 11370
rect 3260 10370 3420 11260
rect 3490 10270 3580 11290
rect 3650 10300 3710 11190
rect 3050 10190 3240 10270
rect 3440 10190 3630 10270
rect 3660 10160 3710 10300
rect 2970 10150 3110 10160
rect 2970 10000 2980 10150
rect 3100 10000 3110 10150
rect 2970 9550 3110 10000
rect 3570 10150 3710 10160
rect 3570 10000 3580 10150
rect 3700 10000 3710 10150
rect 3570 9550 3710 10000
rect 3750 10300 3810 11190
rect 3750 10160 3790 10300
rect 3880 10270 3970 11290
rect 4050 11260 4180 11400
rect 4260 11370 4350 11410
rect 4650 11720 4740 11730
rect 4650 11410 4660 11720
rect 4730 11410 4740 11720
rect 4650 11370 4740 11410
rect 4810 11400 4970 11790
rect 5590 11770 7950 11790
rect 5040 11720 5130 11730
rect 5040 11410 5050 11720
rect 5120 11410 5130 11720
rect 4210 11290 4400 11370
rect 4600 11290 4790 11370
rect 4030 10370 4200 11260
rect 4260 10270 4350 11290
rect 4420 10300 4480 11190
rect 3830 10190 4020 10270
rect 4210 10190 4400 10270
rect 4440 10160 4480 10300
rect 3750 9930 3890 10160
rect 3750 9780 3760 9930
rect 3880 9780 3890 9930
rect 3750 9550 3890 9780
rect 4340 9710 4480 10160
rect 4340 9560 4350 9710
rect 4470 9560 4480 9710
rect 4340 9550 4480 9560
rect 4530 10300 4590 11190
rect 4530 10160 4570 10300
rect 4650 10270 4740 11290
rect 4830 11260 4950 11400
rect 5040 11370 5130 11410
rect 5430 11720 5520 11730
rect 5430 11410 5440 11720
rect 5510 11410 5520 11720
rect 5430 11370 5520 11410
rect 5590 11400 6040 11770
rect 4990 11290 5180 11370
rect 5380 11290 5570 11370
rect 4810 10370 4970 11260
rect 5040 10270 5130 11290
rect 5200 10300 5260 11190
rect 4600 10190 4790 10270
rect 4990 10190 5180 10270
rect 5210 10160 5260 10300
rect 4530 10150 4670 10160
rect 4530 10000 4540 10150
rect 4660 10000 4670 10150
rect 4530 9550 4670 10000
rect 5120 9930 5260 10160
rect 5120 9780 5130 9930
rect 5250 9780 5260 9930
rect 5120 9550 5260 9780
rect 5300 10300 5360 11190
rect 5300 10160 5350 10300
rect 5430 10270 5520 11290
rect 5610 11260 5730 11400
rect 5820 11370 6040 11400
rect 5770 11290 6040 11370
rect 5820 11280 6040 11290
rect 5590 10380 5750 11260
rect 5820 10270 5910 11280
rect 5980 10380 6040 11280
rect 6140 11730 6460 11770
rect 6140 10390 6230 11730
rect 6320 10390 6460 11730
rect 6730 10990 7950 11500
rect 18050 11270 18780 11290
rect 6730 10420 7500 10990
rect 6140 10290 6460 10390
rect 5380 10190 5570 10270
rect 5770 10190 5960 10270
rect 18050 10230 18070 11270
rect 18760 10230 18780 11270
rect 18050 10210 18780 10230
rect 5300 9713 5440 10160
rect 6730 10150 7860 10160
rect 6730 10021 6740 10150
rect 5300 9559 5310 9713
rect 5432 9559 5440 9713
rect 5300 9550 5440 9559
rect 6731 9560 6740 10021
rect 7410 9560 7860 10150
rect 70 9410 5230 9470
rect 70 9320 900 9410
rect 5160 9320 5230 9410
rect 6731 9333 7860 9560
rect 70 9260 5230 9320
rect -812 6892 -582 6930
rect -89 8507 2688 8862
rect -89 8453 0 8507
rect -89 8103 -52 8453
rect -18 8103 0 8453
rect 84 8147 505 8507
rect 1883 8147 2304 8507
rect 2393 8465 2688 8507
rect 2393 8453 7220 8465
rect -89 7945 0 8103
rect 2393 8103 2406 8453
rect 2440 8103 7220 8453
rect 2393 8008 7220 8103
rect -89 7595 -52 7945
rect -18 7595 0 7945
rect -89 7437 0 7595
rect -89 7087 -52 7437
rect -18 7087 0 7437
rect 84 7131 506 7901
rect 1915 7894 3936 7901
rect 1915 7646 3486 7894
rect 3923 7646 3936 7894
rect 1915 7639 3936 7646
rect 4550 7840 7220 8008
rect 4550 7790 5440 7840
rect 4550 7537 4890 7790
rect 2394 7440 4890 7537
rect 4924 7480 5440 7790
rect 6765 7484 7186 7840
rect 4924 7440 4940 7480
rect 2394 7437 4940 7440
rect -89 6929 0 7087
rect -89 6817 -52 6929
rect -2710 6754 -52 6817
rect -2710 6720 -2695 6754
rect -2489 6720 -2331 6754
rect -2125 6720 -1967 6754
rect -1761 6720 -1603 6754
rect -1397 6720 -1239 6754
rect -1033 6720 -875 6754
rect -669 6720 -52 6754
rect -2710 6713 -52 6720
rect -2651 6197 -2169 6618
rect -1923 6198 -1441 6619
rect -1195 6197 -713 6618
rect -615 6579 -52 6713
rect -18 6579 0 6929
rect 1883 6623 2304 7393
rect 2394 7087 2406 7437
rect 2440 7260 4940 7437
rect 2440 7087 4890 7260
rect 2394 6929 4890 7087
rect -615 6421 0 6579
rect -615 6071 -52 6421
rect -18 6071 0 6421
rect 2394 6579 2406 6929
rect 2440 6910 4890 6929
rect 4924 6910 4940 7260
rect 7420 7220 7860 9333
rect 2440 6730 4940 6910
rect 2440 6728 4890 6730
rect 2440 6694 3024 6728
rect 3374 6694 3532 6728
rect 3882 6694 4040 6728
rect 4390 6694 4890 6728
rect 2440 6683 4890 6694
rect 2440 6579 2968 6683
rect 2394 6421 2968 6579
rect -615 5913 0 6071
rect -615 5563 -52 5913
rect -18 5563 0 5913
rect -615 5405 0 5563
rect -615 5055 -52 5405
rect -18 5055 0 5405
rect 84 5099 505 5869
rect 1883 5607 2304 6377
rect 2394 6071 2406 6421
rect 2440 6071 2968 6421
rect 3068 6171 3330 6683
rect 4444 6592 4890 6683
rect 4084 6380 4890 6592
rect 4924 6380 4940 6730
rect 5030 6420 5440 7220
rect 6765 6950 7860 7220
rect 4084 6200 4940 6380
rect 4084 6171 4890 6200
rect 2394 5913 2968 6071
rect 2394 5563 2406 5913
rect 2440 5563 2968 5913
rect 2394 5467 2968 5563
rect 1915 5357 2703 5361
rect 1915 5106 2516 5357
rect 2697 5106 2703 5357
rect 1915 5099 2703 5106
rect -615 4897 0 5055
rect -615 4547 -52 4897
rect -18 4547 0 4897
rect 2395 4897 2688 4994
rect -615 4490 0 4547
rect 84 4490 505 4853
rect 1883 4490 2304 4853
rect 2395 4547 2406 4897
rect 2440 4547 2688 4897
rect 2395 4490 2688 4547
rect -615 4219 2688 4490
rect 2750 4790 2968 5467
rect 4443 5850 4890 6171
rect 4924 5850 4940 6200
rect 4443 5670 4940 5850
rect 4443 5320 4890 5670
rect 4924 5320 4940 5670
rect 5030 5360 5440 6160
rect 6765 5894 7186 6686
rect 4443 5140 4940 5320
rect 4443 4790 4890 5140
rect 4924 4790 4940 5140
rect 2750 4270 3400 4790
rect 2750 4236 3024 4270
rect 3374 4236 3400 4270
rect -615 4080 1780 4219
rect 2750 4200 3400 4236
rect 3480 4140 3930 4790
rect 1810 4130 2080 4140
rect -615 527 394 4080
rect 491 3810 1780 3951
rect 491 527 670 3810
rect 1760 3750 1780 3810
rect 720 3730 1780 3750
rect 1810 3900 1820 4130
rect 2070 3900 2080 4130
rect 720 2670 740 3730
rect 1260 2928 1780 3220
rect 720 2650 1120 2670
rect 1090 2420 1120 2650
rect 720 2400 1120 2420
rect 720 1380 740 2400
rect 720 1360 1120 1380
rect 1090 1130 1120 1360
rect -3015 -2 -2533 419
rect -2286 -2 -1804 419
rect -1559 -1 -1077 420
rect -831 -95 -713 419
rect -615 -40 670 527
rect 720 1110 1120 1130
rect 720 40 740 1110
rect 1260 849 1600 2928
rect 1810 2110 2080 3900
rect 3100 3890 3930 4140
rect 4010 4610 4940 4790
rect 4010 4270 4890 4610
rect 4010 4236 4040 4270
rect 4390 4260 4890 4270
rect 4924 4260 4940 4610
rect 5030 4300 5440 5100
rect 6765 4834 7186 5626
rect 4390 4236 4940 4260
rect 4010 4080 4940 4236
rect 2110 3810 3070 3820
rect 2110 3750 2130 3810
rect 3050 3750 3070 3810
rect 2110 3730 3070 3750
rect 3100 3220 3370 3890
rect 4010 3820 4890 4080
rect 3400 3810 4890 3820
rect 3400 3750 3420 3810
rect 3400 3730 4450 3750
rect 2110 2927 3930 3220
rect 2230 2650 3440 2670
rect 2230 2420 2250 2650
rect 3420 2420 3440 2650
rect 2230 2400 3120 2420
rect 1810 1660 2810 2110
rect 3100 1380 3120 2400
rect 1750 1360 3120 1380
rect 3350 2400 3440 2420
rect 3350 1380 3370 2400
rect 3350 1360 3440 1380
rect 1750 1130 1770 1360
rect 3420 1130 3440 1360
rect 1750 1110 3440 1130
rect 3580 849 3930 2927
rect 4430 2670 4450 3730
rect 4060 2650 4450 2670
rect 4500 3730 4890 3810
rect 4924 3730 4940 4080
rect 4500 3550 4940 3730
rect 4500 3200 4890 3550
rect 4924 3200 4940 3550
rect 5030 3240 5440 4040
rect 6765 3774 7186 4566
rect 4500 3020 4940 3200
rect 4500 2670 4890 3020
rect 4924 2670 4940 3020
rect 4060 2420 4080 2650
rect 4500 2490 4940 2670
rect 4060 2400 4450 2420
rect 4430 1380 4450 2400
rect 4060 1360 4450 1380
rect 4500 2140 4890 2490
rect 4924 2140 4940 2490
rect 5030 2180 5440 2980
rect 6765 2714 7186 3506
rect 6765 2180 7870 2450
rect 4500 1960 4940 2140
rect 4500 1610 4890 1960
rect 4924 1610 4940 1960
rect 4500 1480 4940 1610
rect 5020 1480 5440 1920
rect 6765 1480 7186 1920
rect 4060 1130 4080 1360
rect 4500 1160 7186 1480
rect 4060 1110 4450 1130
rect 1260 560 3930 849
rect 1810 420 2080 440
rect 1810 40 1830 420
rect 720 20 1830 40
rect 2060 40 2080 420
rect 3100 420 3370 440
rect 3100 40 3120 420
rect 2060 20 3120 40
rect 3350 40 3370 420
rect 4430 40 4450 1110
rect 3350 20 4450 40
rect 4500 120 5010 1160
rect 6100 920 7186 1160
rect 7400 850 7870 2180
rect 5230 440 7870 850
rect 6100 120 7970 360
rect 4500 -40 7970 120
rect -615 -95 7970 -40
rect -3701 -104 7970 -95
rect -3701 -138 -3059 -104
rect -2853 -138 -2695 -104
rect -2489 -138 -2331 -104
rect -2125 -138 -1967 -104
rect -1761 -138 -1603 -104
rect -1397 -138 -1239 -104
rect -1033 -138 -875 -104
rect -669 -138 7970 -104
rect -3701 -230 7970 -138
rect -3701 -890 7980 -230
<< via1 >>
rect -2962 11277 -2892 11387
rect -2712 11277 -2632 11387
rect -2322 11277 -2242 11387
rect -1942 11277 -1862 11387
rect -1552 11277 -1472 11387
rect -1162 11277 -1082 11387
rect 1170 11410 1240 11720
rect 1560 11410 1630 11720
rect 1950 11410 2020 11720
rect 1250 9560 1370 9710
rect 2330 11410 2400 11720
rect 2720 11410 2790 11720
rect 1430 9780 1550 9930
rect 2020 10000 2140 10150
rect 3110 11410 3180 11720
rect 3500 11410 3570 11720
rect 2210 9560 2330 9710
rect 2800 9780 2920 9930
rect 3890 11410 3960 11720
rect 4270 11410 4340 11720
rect 2980 10000 3100 10150
rect 3580 10000 3700 10150
rect 4660 11410 4730 11720
rect 5050 11410 5120 11720
rect 3760 9780 3880 9930
rect 4350 9560 4470 9710
rect 5440 11410 5510 11720
rect 4540 10000 4660 10150
rect 5130 9780 5250 9930
rect 13350 11100 18050 11290
rect 18070 10230 18760 11270
rect 5310 9559 5432 9713
rect 6740 9560 7410 10150
rect 3486 7646 3923 7894
rect 103 6636 487 6873
rect 102 6127 487 6367
rect 3589 6190 3825 6573
rect 2516 5106 2697 5357
rect 670 3800 1760 3810
rect 670 3750 1760 3800
rect 1820 3900 2070 4130
rect 670 2420 1090 2650
rect 670 1130 1090 1360
rect 2130 3800 3050 3810
rect 2130 3750 3050 3800
rect 3420 3800 4500 3810
rect 3420 3750 4500 3800
rect 2250 2420 3420 2650
rect 1770 1130 3420 1360
rect 4080 2420 4500 2650
rect 4080 1130 4500 1360
rect 670 -20 4500 20
rect 670 -40 4500 -20
<< metal2 >>
rect -2982 12340 18800 12640
rect -2982 11772 5520 12340
rect -2982 11387 -1072 11772
rect 526 11770 5520 11772
rect 1160 11720 5520 11770
rect -2982 11277 -2962 11387
rect -2892 11277 -2712 11387
rect -2632 11277 -2322 11387
rect -2242 11277 -1942 11387
rect -1862 11277 -1552 11387
rect -1472 11277 -1162 11387
rect -1082 11277 -1072 11387
rect -2982 11267 -1072 11277
rect -529 10160 40 11461
rect 1160 11410 1170 11720
rect 1240 11410 1560 11720
rect 1630 11410 1950 11720
rect 2020 11410 2330 11720
rect 2400 11410 2720 11720
rect 2790 11410 3110 11720
rect 3180 11410 3500 11720
rect 3570 11410 3890 11720
rect 3960 11410 4270 11720
rect 4340 11410 4660 11720
rect 4730 11410 5050 11720
rect 5120 11410 5440 11720
rect 5510 11410 5520 11720
rect 1160 11400 5520 11410
rect 13330 11290 18800 12340
rect 13330 11100 13350 11290
rect 18050 11270 18800 11290
rect 18050 11100 18070 11270
rect 13330 11080 18070 11100
rect -529 10150 7420 10160
rect -529 10000 2020 10150
rect 2140 10000 2980 10150
rect 3100 10000 3580 10150
rect 3700 10000 4540 10150
rect 4660 10010 6740 10150
rect 4660 10000 5440 10010
rect -529 9990 5440 10000
rect 620 9940 1259 9941
rect 620 9930 5681 9940
rect 620 9780 1430 9930
rect 1550 9780 2800 9930
rect 2920 9780 3760 9930
rect 3880 9780 5130 9930
rect 5250 9780 5681 9930
rect 620 9770 5681 9780
rect 620 9224 1057 9770
rect 1230 9713 5681 9720
rect 1230 9710 5310 9713
rect 1230 9560 1250 9710
rect 1370 9560 2210 9710
rect 2330 9560 4350 9710
rect 4470 9560 5310 9710
rect 1230 9559 5310 9560
rect 5432 9559 5681 9713
rect 1230 9550 5681 9559
rect 5756 9560 6740 10010
rect 7410 9560 7420 10150
rect 5756 9551 7420 9560
rect 6731 9550 7420 9551
rect -506 8917 1057 9224
rect -506 6378 -322 8917
rect 1595 8867 1981 9550
rect 7650 9232 8490 10270
rect 18030 10230 18070 11080
rect 18760 10230 18800 11270
rect 18030 10190 18800 10230
rect 6030 9230 8490 9232
rect -262 8625 1981 8867
rect 2509 8790 8490 9230
rect -262 6885 -15 8625
rect 2509 8243 2858 8790
rect -262 6873 505 6885
rect -262 6636 103 6873
rect 487 6636 505 6873
rect -262 6623 505 6636
rect -506 6367 505 6378
rect -506 6127 102 6367
rect 487 6127 505 6367
rect -506 6115 505 6127
rect 2509 5368 2859 8243
rect 3480 8130 7880 8670
rect 3480 7894 3930 8130
rect 3480 7646 3486 7894
rect 3923 7646 3930 7894
rect 3480 6573 3930 7646
rect 3480 6190 3589 6573
rect 3825 6190 3930 6573
rect 3480 6171 3930 6190
rect 2509 5357 2860 5368
rect 2509 5106 2516 5357
rect 2697 5106 2860 5357
rect 2509 4140 2860 5106
rect 1810 4130 2860 4140
rect 1810 3900 1820 4130
rect 2070 3900 2860 4130
rect 1810 3890 2860 3900
rect 630 3810 4550 3840
rect 630 3750 670 3810
rect 1760 3750 2130 3810
rect 3050 3750 3420 3810
rect 4500 3750 4550 3810
rect 630 3730 4550 3750
rect 630 2650 4540 2670
rect 630 2420 670 2650
rect 1090 2420 2250 2650
rect 3420 2420 4080 2650
rect 4500 2420 4540 2650
rect 630 2400 4540 2420
rect 630 1360 4550 1380
rect 630 1130 670 1360
rect 1090 1130 1770 1360
rect 3420 1130 4080 1360
rect 4500 1130 4550 1360
rect 630 1110 4550 1130
rect 630 20 4550 40
rect 630 -40 670 20
rect 4500 -40 4550 20
rect 630 -60 4550 -40
use bmbgota  bmbgota_0
timestamp 1725107840
transform 1 0 9631 0 1 8620
box -1820 -9510 9170 3660
use sky130_fd_pr__pfet_g5v0d10v5_SSAD3V  sky130_fd_pr__pfet_g5v0d10v5_SSAD3V_0
timestamp 1725192216
transform -1 0 -3012 0 -1 9144
box -174 -2100 174 2100
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_0
timestamp 1646940291
transform 1 0 818 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_1
timestamp 1646940291
transform 1 0 1206 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_2
timestamp 1646940291
transform 1 0 1594 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_3
timestamp 1646940291
transform 1 0 1982 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_4
timestamp 1646940291
transform 1 0 2370 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_5
timestamp 1646940291
transform 1 0 2758 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_6
timestamp 1646940291
transform 1 0 3146 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_7
timestamp 1646940291
transform 1 0 3534 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_8
timestamp 1646940291
transform 1 0 3922 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_9
timestamp 1646940291
transform 1 0 4310 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_10
timestamp 1646940291
transform 1 0 4698 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_11
timestamp 1646940291
transform 1 0 5086 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_12
timestamp 1646940291
transform 1 0 5474 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_XYTFBH  sky130_fd_pr__pfet_g5v0d10v5_XYTFBH_13
timestamp 1646940291
transform 1 0 5862 0 1 10781
box -224 -600 224 600
use sky130_fd_pr__pfet_g5v0d10v5_ZL3LRV  sky130_fd_pr__pfet_g5v0d10v5_ZL3LRV_0
timestamp 1646941581
transform -1 0 -1121 0 -1 9144
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_ZL3LRV  sky130_fd_pr__pfet_g5v0d10v5_ZL3LRV_1
timestamp 1646941581
transform -1 0 -1509 0 -1 9144
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_ZL3LRV  sky130_fd_pr__pfet_g5v0d10v5_ZL3LRV_2
timestamp 1646941581
transform -1 0 -1897 0 -1 9144
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_ZL3LRV  sky130_fd_pr__pfet_g5v0d10v5_ZL3LRV_3
timestamp 1646941581
transform -1 0 -2285 0 -1 9144
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_ZL3LRV  sky130_fd_pr__pfet_g5v0d10v5_ZL3LRV_4
timestamp 1646941581
transform -1 0 -2673 0 -1 9144
box -224 -2100 224 2100
use sky130_fd_pr__res_xhigh_po_0p69_7V2R7J  sky130_fd_pr__res_xhigh_po_0p69_7V2R7J_0
timestamp 1724871964
transform 1 0 -2228 0 1 3308
box -235 -3482 235 3482
use sky130_fd_pr__res_xhigh_po_0p69_7V2R7J  sky130_fd_pr__res_xhigh_po_0p69_7V2R7J_1
timestamp 1724871964
transform 1 0 -2956 0 1 3308
box -235 -3482 235 3482
use sky130_fd_pr__res_xhigh_po_0p69_7V2R7J  sky130_fd_pr__res_xhigh_po_0p69_7V2R7J_2
timestamp 1724871964
transform 1 0 -772 0 1 3308
box -235 -3482 235 3482
use sky130_fd_pr__res_xhigh_po_0p69_7V2R7J  sky130_fd_pr__res_xhigh_po_0p69_7V2R7J_3
timestamp 1724871964
transform 1 0 -1864 0 1 3308
box -235 -3482 235 3482
use sky130_fd_pr__res_xhigh_po_0p69_7V2R7J  sky130_fd_pr__res_xhigh_po_0p69_7V2R7J_4
timestamp 1724871964
transform 1 0 -1500 0 1 3308
box -235 -3482 235 3482
use sky130_fd_pr__res_xhigh_po_0p69_7V2R7J  sky130_fd_pr__res_xhigh_po_0p69_7V2R7J_5
timestamp 1724871964
transform 1 0 -1136 0 1 3308
box -235 -3482 235 3482
use sky130_fd_pr__res_xhigh_po_0p69_7V2R7J  sky130_fd_pr__res_xhigh_po_0p69_7V2R7J_6
timestamp 1724871964
transform 1 0 -2592 0 1 3308
box -235 -3482 235 3482
use sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8  sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8_0
timestamp 1725102575
transform 0 1 1194 -1 0 4722
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8  sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8_1
timestamp 1725102575
transform 0 1 1194 -1 0 8278
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8  sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8_2
timestamp 1725102575
transform 0 1 1194 -1 0 7770
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8  sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8_3
timestamp 1725102575
transform 0 1 1194 -1 0 7262
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8  sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8_4
timestamp 1725102575
transform 0 1 1194 -1 0 6754
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8  sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8_5
timestamp 1725102575
transform 0 1 1194 -1 0 6246
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8  sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8_6
timestamp 1725102575
transform 0 1 1194 -1 0 5738
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8  sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8_7
timestamp 1725102575
transform 0 1 1194 -1 0 5230
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8  sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8_8
timestamp 1725102575
transform 1 0 4215 0 1 5482
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8  sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8_9
timestamp 1725102575
transform 1 0 3199 0 1 5482
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8  sky130_fd_pr__res_xhigh_po_1p41_2SU5Y8_10
timestamp 1725102575
transform 1 0 3707 0 1 5482
box -307 -1282 307 1282
use sky130_fd_pr__res_xhigh_po_1p41_T77NL5  sky130_fd_pr__res_xhigh_po_1p41_T77NL5_0
timestamp 1725107131
transform 0 1 6106 -1 0 7615
box -307 -1252 307 1252
use sky130_fd_pr__res_xhigh_po_1p41_T77NL5  sky130_fd_pr__res_xhigh_po_1p41_T77NL5_1
timestamp 1725107131
transform 0 1 6106 -1 0 1785
box -307 -1252 307 1252
use sky130_fd_pr__res_xhigh_po_1p41_T77NL5  sky130_fd_pr__res_xhigh_po_1p41_T77NL5_2
timestamp 1725107131
transform 0 1 6106 -1 0 7085
box -307 -1252 307 1252
use sky130_fd_pr__res_xhigh_po_1p41_T77NL5  sky130_fd_pr__res_xhigh_po_1p41_T77NL5_3
timestamp 1725107131
transform 0 1 6106 -1 0 6555
box -307 -1252 307 1252
use sky130_fd_pr__res_xhigh_po_1p41_T77NL5  sky130_fd_pr__res_xhigh_po_1p41_T77NL5_4
timestamp 1725107131
transform 0 1 6106 -1 0 6025
box -307 -1252 307 1252
use sky130_fd_pr__res_xhigh_po_1p41_T77NL5  sky130_fd_pr__res_xhigh_po_1p41_T77NL5_5
timestamp 1725107131
transform 0 1 6106 -1 0 5495
box -307 -1252 307 1252
use sky130_fd_pr__res_xhigh_po_1p41_T77NL5  sky130_fd_pr__res_xhigh_po_1p41_T77NL5_6
timestamp 1725107131
transform 0 1 6106 -1 0 4965
box -307 -1252 307 1252
use sky130_fd_pr__res_xhigh_po_1p41_T77NL5  sky130_fd_pr__res_xhigh_po_1p41_T77NL5_7
timestamp 1725107131
transform 0 1 6106 -1 0 4435
box -307 -1252 307 1252
use sky130_fd_pr__res_xhigh_po_1p41_T77NL5  sky130_fd_pr__res_xhigh_po_1p41_T77NL5_8
timestamp 1725107131
transform 0 1 6106 -1 0 3905
box -307 -1252 307 1252
use sky130_fd_pr__res_xhigh_po_1p41_T77NL5  sky130_fd_pr__res_xhigh_po_1p41_T77NL5_9
timestamp 1725107131
transform 0 1 6106 -1 0 3375
box -307 -1252 307 1252
use sky130_fd_pr__res_xhigh_po_1p41_T77NL5  sky130_fd_pr__res_xhigh_po_1p41_T77NL5_10
timestamp 1725107131
transform 0 1 6106 -1 0 2845
box -307 -1252 307 1252
use sky130_fd_pr__res_xhigh_po_1p41_T77NL5  sky130_fd_pr__res_xhigh_po_1p41_T77NL5_11
timestamp 1725107131
transform 0 1 6106 -1 0 2315
box -307 -1252 307 1252
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 630 0 1 -70
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 1918 0 1 -70
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 3206 0 1 -70
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 630 0 1 1218
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 1918 0 1 1218
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 3206 0 1 1218
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 630 0 1 2506
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1723858470
transform 1 0 1918 0 1 2506
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1723858470
transform 1 0 3206 0 1 2506
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9
timestamp 1723858470
transform 1 0 4855 0 1 -29
box 0 0 1340 1340
<< labels >>
flabel metal1 6730 10420 7500 10990 0 FreeSans 1600 0 0 0 IB
port 2 nsew
flabel metal2 -512 10013 19 11443 0 FreeSans 1600 0 0 0 VREF
port 3 nsew
flabel metal1 -3694 -883 -3534 -13 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal1 -3681 11680 -3521 12550 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
<< end >>
