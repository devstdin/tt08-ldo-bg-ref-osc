magic
tech sky130A
magscale 1 2
timestamp 1725466509
<< metal1 >>
rect 27207 44829 27350 44836
rect 27207 44700 27214 44829
rect 27343 44700 27350 44829
rect 27207 44693 27350 44700
rect 800 44132 1200 44152
rect 800 33214 820 44132
rect 1180 42958 1200 44132
rect 1419 44118 2945 44323
rect 1419 43176 1433 44118
rect 1765 43176 2945 44118
rect 1419 43161 2945 43176
rect 1180 40079 2723 42958
rect 1180 39751 1200 40079
rect 1180 33214 1860 39751
rect 24192 38726 25295 38806
rect 24192 38009 24371 38726
rect 24437 38009 25295 38726
rect 24192 37751 25295 38009
rect 24192 34648 24369 37751
rect 24191 34196 24369 34648
rect 800 33194 1860 33214
rect 931 33035 1860 33194
rect 24192 33341 24369 34196
rect 24439 33341 25295 37751
rect 24192 33212 25295 33341
rect 24192 33203 27129 33212
rect 16199 33035 16590 33154
rect 24192 33035 26674 33203
rect 931 32713 26674 33035
rect 27118 32713 27129 33203
rect 931 32702 27129 32713
rect 931 32701 25295 32702
rect 27214 32529 27343 44693
rect 27649 44602 27793 44609
rect 27649 44473 27656 44602
rect 27785 44473 27793 44602
rect 27649 44465 27793 44473
rect 800 32401 1200 32421
rect 800 1020 820 32401
rect 1180 26543 1200 32401
rect 1401 32387 2052 32419
rect 1401 31221 1432 32387
rect 1765 31221 2052 32387
rect 25628 32400 27343 32529
rect 25628 31749 25757 32400
rect 27656 32288 27785 44465
rect 28120 44273 28264 44280
rect 28120 44144 28127 44273
rect 28256 44144 28264 44273
rect 28120 44137 28264 44144
rect 25836 32159 27785 32288
rect 25836 31749 25965 32159
rect 28127 32060 28256 44137
rect 26154 31931 28256 32060
rect 26154 31748 26283 31931
rect 1401 31206 2052 31221
rect 12297 31421 13067 31443
rect 12297 30221 12319 31421
rect 13045 30221 13067 31421
rect 12297 30199 13067 30221
rect 1180 18888 1918 26543
rect 27740 26286 27967 26537
rect 27740 26124 27746 26286
rect 27961 26124 27967 26286
rect 27740 26118 27967 26124
rect 1180 9244 1200 18888
rect 1409 18750 5261 18764
rect 1409 15080 1432 18750
rect 1764 15080 5261 18750
rect 1409 15066 5261 15080
rect 3908 14104 5066 14124
rect 3908 13444 3927 14104
rect 4704 13444 5066 14104
rect 3908 13424 5066 13444
rect 3983 10303 5434 10313
rect 3983 9623 3992 10303
rect 4404 9623 5434 10303
rect 3983 9615 5434 9623
rect 1180 7843 5430 9244
rect 1180 1020 1200 7843
rect 3983 3412 5394 3424
rect 3983 2806 3995 3412
rect 4402 2806 5394 3412
rect 3983 2794 5394 2806
rect 800 1000 1200 1020
<< via1 >>
rect 27214 44700 27343 44829
rect 820 33214 1180 44132
rect 1433 43176 1765 44118
rect 26674 32713 27118 33203
rect 27656 44473 27785 44602
rect 820 1020 1180 32401
rect 1432 31221 1765 32387
rect 28127 44144 28256 44273
rect 12319 30221 13045 31421
rect 27746 26124 27961 26286
rect 1432 15080 1764 18750
rect 3927 13444 4704 14104
rect 3992 9623 4404 10303
rect 3995 2806 4402 3412
<< metal2 >>
rect 25815 44701 25824 44830
rect 25953 44829 25962 44830
rect 27207 44829 27350 44836
rect 25953 44701 27214 44829
rect 25824 44700 27214 44701
rect 27343 44700 27350 44829
rect 27207 44693 27350 44700
rect 27649 44602 27793 44609
rect 26158 44473 26167 44602
rect 26296 44473 27656 44602
rect 27785 44473 27793 44602
rect 27649 44465 27793 44473
rect 28120 44273 28264 44280
rect 800 44132 1200 44152
rect 800 33214 820 44132
rect 1180 33214 1200 44132
rect 800 33194 1200 33214
rect 1400 44132 1800 44152
rect 16846 44144 16855 44273
rect 16984 44144 28127 44273
rect 28256 44144 28264 44273
rect 28120 44137 28264 44144
rect 1400 33214 1420 44132
rect 1780 33214 1800 44132
rect 26395 38883 28859 39017
rect 25507 38843 28859 38883
rect 1400 33194 1800 33214
rect 26663 33203 27129 33212
rect 26663 32713 26674 33203
rect 27118 32713 27129 33203
rect 800 32401 1200 32421
rect 800 1020 820 32401
rect 1180 1020 1200 32401
rect 800 1000 1200 1020
rect 1400 32401 1800 32421
rect 1400 1020 1420 32401
rect 1780 1020 1800 32401
rect 26663 31749 27129 32713
rect 28067 33026 28516 33043
rect 28067 32595 28078 33026
rect 28506 32595 28516 33026
rect 28067 32093 28516 32595
rect 28067 31747 28517 32093
rect 12297 31421 13067 31443
rect 12297 30221 12319 31421
rect 13045 30221 13067 31421
rect 12297 30199 13067 30221
rect 28685 26292 28859 38843
rect 27735 26286 28859 26292
rect 27735 26124 27746 26286
rect 27961 26124 28859 26286
rect 27735 26118 28859 26124
rect 3907 14104 4724 14124
rect 3907 13444 3927 14104
rect 4704 13444 4724 14104
rect 3907 13424 4724 13444
rect 3983 10303 4414 10313
rect 3983 9623 3992 10303
rect 4404 9623 4414 10303
rect 3983 3412 4414 9623
rect 23886 7974 24952 7984
rect 23886 6885 24428 7974
rect 24939 6885 24952 7974
rect 23886 6874 24952 6885
rect 3983 2806 3995 3412
rect 4402 2806 4414 3412
rect 3983 2794 4414 2806
rect 1400 1000 1800 1020
<< via2 >>
rect 25824 44701 25953 44830
rect 26167 44473 26296 44602
rect 820 33214 1180 44132
rect 16855 44144 16984 44273
rect 1420 44118 1780 44132
rect 1420 43176 1433 44118
rect 1433 43176 1765 44118
rect 1765 43176 1780 44118
rect 1420 33214 1780 43176
rect 21820 38758 22592 39034
rect 23002 38849 23870 39122
rect 820 1020 1180 32401
rect 1420 32387 1780 32401
rect 1420 31221 1432 32387
rect 1432 31221 1765 32387
rect 1765 31221 1780 32387
rect 1420 18750 1780 31221
rect 1420 15080 1432 18750
rect 1432 15080 1764 18750
rect 1764 15080 1780 18750
rect 1420 1020 1780 15080
rect 28078 32595 28506 33026
rect 5055 29792 5586 31222
rect 12319 30221 13045 31421
rect 3927 13444 4704 14104
rect 24428 6885 24939 7974
rect 4790 3715 5234 4550
<< metal3 >>
rect 25819 44830 25958 44835
rect 23943 44701 23949 44830
rect 24078 44701 25824 44830
rect 25953 44701 25958 44830
rect 25819 44696 25958 44701
rect 26162 44602 26301 44607
rect 24497 44473 24503 44602
rect 24632 44473 26167 44602
rect 26296 44473 26301 44602
rect 26162 44468 26301 44473
rect 16850 44273 16989 44278
rect 800 44132 1200 44152
rect 800 33214 820 44132
rect 1180 33214 1200 44132
rect 800 33194 1200 33214
rect 1400 44132 1800 44152
rect 15664 44144 15670 44273
rect 15799 44144 16855 44273
rect 16984 44144 16989 44273
rect 16850 44139 16989 44144
rect 1400 33214 1420 44132
rect 1780 33214 1800 44132
rect 2544 41343 23882 41360
rect 2544 40487 2557 41343
rect 3328 40487 23882 41343
rect 2544 40472 23882 40487
rect 12283 39970 22605 40003
rect 12283 39222 12316 39970
rect 13047 39222 22605 39970
rect 12283 39204 22605 39222
rect 21806 39034 22605 39204
rect 21806 38758 21820 39034
rect 22592 38758 22605 39034
rect 22994 39122 23882 40472
rect 22994 38849 23002 39122
rect 23870 38849 23882 39122
rect 22994 38840 23882 38849
rect 21806 38745 22605 38758
rect 1400 33194 1800 33214
rect 202 33027 28524 33036
rect 202 32594 210 33027
rect 592 33026 28524 33027
rect 592 32595 28078 33026
rect 28506 32595 28524 33026
rect 592 32594 28524 32595
rect 202 32584 28524 32594
rect 800 32401 1200 32421
rect 800 1020 820 32401
rect 1180 1020 1200 32401
rect 800 1000 1200 1020
rect 1400 32401 1800 32421
rect 1400 1020 1420 32401
rect 1780 1020 1800 32401
rect 12297 31421 13067 31443
rect 5038 31222 5607 31240
rect 5038 29792 5055 31222
rect 5586 29792 5607 31222
rect 12297 30221 12319 31421
rect 13045 30221 13067 31421
rect 12297 30199 13067 30221
rect 5038 29769 5607 29792
rect 3907 14104 4724 14124
rect 3907 13444 3927 14104
rect 4704 13444 4724 14104
rect 3907 13424 4724 13444
rect 24416 7974 27412 7984
rect 24416 6885 24428 7974
rect 24939 7972 27412 7974
rect 24939 6886 26848 7972
rect 27401 6886 27412 7972
rect 24939 6885 27412 6886
rect 24416 6874 27412 6885
rect 2545 4551 5250 4564
rect 2545 3716 2558 4551
rect 3333 4550 5250 4551
rect 3333 3716 4790 4550
rect 2545 3715 4790 3716
rect 5234 3715 5250 4550
rect 2545 3704 5250 3715
rect 1400 1000 1800 1020
<< via3 >>
rect 23949 44701 24078 44830
rect 24503 44473 24632 44602
rect 820 33214 1180 44132
rect 15670 44144 15799 44273
rect 1420 33214 1780 44132
rect 2557 40487 3328 41343
rect 12316 39222 13047 39970
rect 210 32594 592 33027
rect 820 1020 1180 32401
rect 1420 1020 1780 32401
rect 5055 29792 5586 31222
rect 12319 30221 13045 31421
rect 3927 13444 4704 14104
rect 26848 6886 27401 7972
rect 2558 3716 3333 4551
<< metal4 >>
rect 3006 44969 3066 45152
rect 3558 44969 3618 45152
rect 4110 44969 4170 45152
rect 4662 44969 4722 45152
rect 5214 44969 5274 45152
rect 5766 44969 5826 45152
rect 6318 44969 6378 45152
rect 6870 44969 6930 45152
rect 7422 44969 7482 45152
rect 7974 44969 8034 45152
rect 8526 44969 8586 45152
rect 9078 44969 9138 45152
rect 9630 44969 9690 45152
rect 10182 44969 10242 45152
rect 10734 44969 10794 45152
rect 11286 44969 11346 45152
rect 11838 44969 11898 45152
rect 12390 44969 12450 45152
rect 12942 44969 13002 45152
rect 13494 44969 13554 45152
rect 14046 44969 14106 45152
rect 14598 44969 14658 45152
rect 15150 44969 15210 45152
rect 15702 44974 15762 45152
rect 912 44784 15210 44969
rect 912 44152 1097 44784
rect 15670 44274 15799 44974
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44968 24042 45152
rect 23949 44831 24078 44968
rect 24534 44966 24594 45152
rect 23948 44830 24079 44831
rect 23948 44701 23949 44830
rect 24078 44701 24079 44830
rect 23948 44700 24079 44701
rect 24503 44603 24632 44966
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 24502 44602 24633 44603
rect 24502 44473 24503 44602
rect 24632 44473 24633 44602
rect 24502 44472 24633 44473
rect 15669 44273 15800 44274
rect 200 33027 600 44152
rect 200 32594 210 33027
rect 592 32594 600 33027
rect 200 1000 600 32594
rect 800 44132 1200 44152
rect 800 33214 820 44132
rect 1180 33214 1200 44132
rect 800 32401 1200 33214
rect 800 1020 820 32401
rect 1180 1020 1200 32401
rect 800 1000 1200 1020
rect 1400 44132 1800 44152
rect 15669 44144 15670 44273
rect 15799 44144 15800 44273
rect 15669 44143 15800 44144
rect 1400 33214 1420 44132
rect 1780 33214 1800 44132
rect 1400 32401 1800 33214
rect 1400 1020 1420 32401
rect 1780 1020 1800 32401
rect 2545 41343 3350 41360
rect 2545 40487 2557 41343
rect 3328 40487 3350 41343
rect 2545 4551 3350 40487
rect 12297 39970 13067 39987
rect 12297 39222 12316 39970
rect 13047 39222 13067 39970
rect 12297 31421 13067 39222
rect 3907 31222 5607 31240
rect 3907 29792 5055 31222
rect 5586 29792 5607 31222
rect 12297 30221 12319 31421
rect 13045 30221 13067 31421
rect 12297 30199 13067 30221
rect 3907 29769 5607 29792
rect 3907 14104 4724 29769
rect 3907 13444 3927 14104
rect 4704 13444 4724 14104
rect 3907 13424 4724 13444
rect 2545 3716 2558 4551
rect 3333 3716 3350 4551
rect 2545 3704 3350 3716
rect 26836 7972 27414 7984
rect 26836 6886 26848 7972
rect 27401 6886 27414 7972
rect 1400 1000 1800 1020
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 26836 170 27414 6886
rect 27234 0 27414 170
use bmbg  bmbg_0 ../ip/bmbg/magic
timestamp 1725192368
transform 1 0 5567 0 1 19779
box -3701 -890 18801 12640
use ldo  ldo_0 ../ip/ldo/magic
timestamp 1725202063
transform 1 0 3188 0 1 8444
box 1590 -7310 21171 10320
use riosc  riosc_0 ../ip/riosc/magic
timestamp 1725202727
transform 0 1 25155 -1 0 30629
box -1218 259 4183 3362
use vthref  vthref_0 ../ip/vthref_tt/magic
timestamp 1725184256
transform 1 0 7516 0 1 39413
box -5663 -6320 16868 4909
use vthref_source  vthref_source_0 ../ip/vthref_tt/magic
timestamp 1724418000
transform 1 0 10029 0 1 39416
box 14026 -573 16868 4906
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1400 1000 1800 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
