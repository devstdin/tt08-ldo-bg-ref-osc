magic
tech sky130A
magscale 1 2
timestamp 1725107131
<< pwell >>
rect -307 -1252 307 1252
<< psubdiff >>
rect -271 1182 -175 1216
rect 175 1182 271 1216
rect -271 -1182 -237 1182
rect 237 -1182 271 1182
rect -271 -1216 -175 -1182
rect 175 -1216 271 -1182
<< psubdiffcont >>
rect -175 1182 175 1216
rect -175 -1216 175 -1182
<< xpolycontact >>
rect -141 654 141 1086
rect -141 -1086 141 -654
<< xpolyres >>
rect -141 -654 141 654
<< locali >>
rect -271 1182 -175 1216
rect 175 1182 271 1216
rect -271 -1182 -237 1182
rect 237 -1182 271 1182
rect -271 -1216 -175 -1182
rect 175 -1216 271 -1182
<< viali >>
rect -125 671 125 1068
rect -125 -1068 125 -671
<< metal1 >>
rect -131 1068 131 1080
rect -131 671 -125 1068
rect 125 671 131 1068
rect -131 659 131 671
rect -131 -671 131 -659
rect -131 -1068 -125 -671
rect 125 -1068 131 -671
rect -131 -1080 131 -1068
<< properties >>
string FIXED_BBOX -254 -1199 254 1199
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 6.7 m 1 nx 1 wmin 1.410 lmin 0.50 class resistor rho 2000 val 9.77k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 0 grc 0 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
