magic
tech sky130A
magscale 1 2
timestamp 1650714605
<< error_p >>
rect -4549 4490 -4329 8550
rect -8628 4350 -4329 4490
rect -4309 4490 -4089 8550
rect -230 4490 -10 8550
rect -4309 4350 -10 4490
rect 10 4490 230 8550
rect 4089 4490 4309 8550
rect 10 4350 4309 4490
rect 4329 4490 4549 8550
rect 4329 4350 8628 4490
rect -8628 4110 -4329 4250
rect -4549 190 -4329 4110
rect -8628 50 -4329 190
rect -4309 4110 -10 4250
rect -4309 190 -4089 4110
rect -230 190 -10 4110
rect -4309 50 -10 190
rect 10 4110 4309 4250
rect 10 190 230 4110
rect 4089 190 4309 4110
rect 10 50 4309 190
rect 4329 4110 8628 4250
rect 4329 190 4549 4110
rect 4329 50 8628 190
rect -8628 -190 -4329 -50
rect -4549 -4110 -4329 -190
rect -8628 -4250 -4329 -4110
rect -4309 -190 -10 -50
rect -4309 -4110 -4089 -190
rect -230 -4110 -10 -190
rect -4309 -4250 -10 -4110
rect 10 -190 4309 -50
rect 10 -4110 230 -190
rect 4089 -4110 4309 -190
rect 10 -4250 4309 -4110
rect 4329 -190 8628 -50
rect 4329 -4110 4549 -190
rect 4329 -4250 8628 -4110
rect -8628 -4490 -4329 -4350
rect -4549 -8550 -4329 -4490
rect -4309 -4490 -10 -4350
rect -4309 -8550 -4089 -4490
rect -230 -8550 -10 -4490
rect 10 -4490 4309 -4350
rect 10 -8550 230 -4490
rect 4089 -8550 4309 -4490
rect 4329 -4490 8628 -4350
rect 4329 -8550 4549 -4490
<< metal3 >>
rect -8628 8522 -4329 8550
rect -8628 4378 -4413 8522
rect -4349 4378 -4329 8522
rect -8628 4350 -4329 4378
rect -4309 8522 -10 8550
rect -4309 4378 -94 8522
rect -30 4378 -10 8522
rect -4309 4350 -10 4378
rect 10 8522 4309 8550
rect 10 4378 4225 8522
rect 4289 4378 4309 8522
rect 10 4350 4309 4378
rect 4329 8522 8628 8550
rect 4329 4378 8544 8522
rect 8608 4378 8628 8522
rect 4329 4350 8628 4378
rect -8628 4222 -4329 4250
rect -8628 78 -4413 4222
rect -4349 78 -4329 4222
rect -8628 50 -4329 78
rect -4309 4222 -10 4250
rect -4309 78 -94 4222
rect -30 78 -10 4222
rect -4309 50 -10 78
rect 10 4222 4309 4250
rect 10 78 4225 4222
rect 4289 78 4309 4222
rect 10 50 4309 78
rect 4329 4222 8628 4250
rect 4329 78 8544 4222
rect 8608 78 8628 4222
rect 4329 50 8628 78
rect -8628 -78 -4329 -50
rect -8628 -4222 -4413 -78
rect -4349 -4222 -4329 -78
rect -8628 -4250 -4329 -4222
rect -4309 -78 -10 -50
rect -4309 -4222 -94 -78
rect -30 -4222 -10 -78
rect -4309 -4250 -10 -4222
rect 10 -78 4309 -50
rect 10 -4222 4225 -78
rect 4289 -4222 4309 -78
rect 10 -4250 4309 -4222
rect 4329 -78 8628 -50
rect 4329 -4222 8544 -78
rect 8608 -4222 8628 -78
rect 4329 -4250 8628 -4222
rect -8628 -4378 -4329 -4350
rect -8628 -8522 -4413 -4378
rect -4349 -8522 -4329 -4378
rect -8628 -8550 -4329 -8522
rect -4309 -4378 -10 -4350
rect -4309 -8522 -94 -4378
rect -30 -8522 -10 -4378
rect -4309 -8550 -10 -8522
rect 10 -4378 4309 -4350
rect 10 -8522 4225 -4378
rect 4289 -8522 4309 -4378
rect 10 -8550 4309 -8522
rect 4329 -4378 8628 -4350
rect 4329 -8522 8544 -4378
rect 8608 -8522 8628 -4378
rect 4329 -8550 8628 -8522
<< via3 >>
rect -4413 4378 -4349 8522
rect -94 4378 -30 8522
rect 4225 4378 4289 8522
rect 8544 4378 8608 8522
rect -4413 78 -4349 4222
rect -94 78 -30 4222
rect 4225 78 4289 4222
rect 8544 78 8608 4222
rect -4413 -4222 -4349 -78
rect -94 -4222 -30 -78
rect 4225 -4222 4289 -78
rect 8544 -4222 8608 -78
rect -4413 -8522 -4349 -4378
rect -94 -8522 -30 -4378
rect 4225 -8522 4289 -4378
rect 8544 -8522 8608 -4378
<< mimcap >>
rect -8528 8410 -4528 8450
rect -8528 4490 -8488 8410
rect -4568 4490 -4528 8410
rect -8528 4450 -4528 4490
rect -4209 8410 -209 8450
rect -4209 4490 -4169 8410
rect -249 4490 -209 8410
rect -4209 4450 -209 4490
rect 110 8410 4110 8450
rect 110 4490 150 8410
rect 4070 4490 4110 8410
rect 110 4450 4110 4490
rect 4429 8410 8429 8450
rect 4429 4490 4469 8410
rect 8389 4490 8429 8410
rect 4429 4450 8429 4490
rect -8528 4110 -4528 4150
rect -8528 190 -8488 4110
rect -4568 190 -4528 4110
rect -8528 150 -4528 190
rect -4209 4110 -209 4150
rect -4209 190 -4169 4110
rect -249 190 -209 4110
rect -4209 150 -209 190
rect 110 4110 4110 4150
rect 110 190 150 4110
rect 4070 190 4110 4110
rect 110 150 4110 190
rect 4429 4110 8429 4150
rect 4429 190 4469 4110
rect 8389 190 8429 4110
rect 4429 150 8429 190
rect -8528 -190 -4528 -150
rect -8528 -4110 -8488 -190
rect -4568 -4110 -4528 -190
rect -8528 -4150 -4528 -4110
rect -4209 -190 -209 -150
rect -4209 -4110 -4169 -190
rect -249 -4110 -209 -190
rect -4209 -4150 -209 -4110
rect 110 -190 4110 -150
rect 110 -4110 150 -190
rect 4070 -4110 4110 -190
rect 110 -4150 4110 -4110
rect 4429 -190 8429 -150
rect 4429 -4110 4469 -190
rect 8389 -4110 8429 -190
rect 4429 -4150 8429 -4110
rect -8528 -4490 -4528 -4450
rect -8528 -8410 -8488 -4490
rect -4568 -8410 -4528 -4490
rect -8528 -8450 -4528 -8410
rect -4209 -4490 -209 -4450
rect -4209 -8410 -4169 -4490
rect -249 -8410 -209 -4490
rect -4209 -8450 -209 -8410
rect 110 -4490 4110 -4450
rect 110 -8410 150 -4490
rect 4070 -8410 4110 -4490
rect 110 -8450 4110 -8410
rect 4429 -4490 8429 -4450
rect 4429 -8410 4469 -4490
rect 8389 -8410 8429 -4490
rect 4429 -8450 8429 -8410
<< mimcapcontact >>
rect -8488 4490 -4568 8410
rect -4169 4490 -249 8410
rect 150 4490 4070 8410
rect 4469 4490 8389 8410
rect -8488 190 -4568 4110
rect -4169 190 -249 4110
rect 150 190 4070 4110
rect 4469 190 8389 4110
rect -8488 -4110 -4568 -190
rect -4169 -4110 -249 -190
rect 150 -4110 4070 -190
rect 4469 -4110 8389 -190
rect -8488 -8410 -4568 -4490
rect -4169 -8410 -249 -4490
rect 150 -8410 4070 -4490
rect 4469 -8410 8389 -4490
<< metal4 >>
rect -6580 8411 -6476 8600
rect -4460 8538 -4356 8600
rect -4460 8522 -4333 8538
rect -8489 8410 -4567 8411
rect -8489 4490 -8488 8410
rect -4568 4490 -4567 8410
rect -8489 4489 -4567 4490
rect -6580 4111 -6476 4489
rect -4460 4378 -4413 8522
rect -4349 4378 -4333 8522
rect -2261 8411 -2157 8600
rect -141 8538 -37 8600
rect -141 8522 -14 8538
rect -4170 8410 -248 8411
rect -4170 4490 -4169 8410
rect -249 4490 -248 8410
rect -4170 4489 -248 4490
rect -4460 4362 -4333 4378
rect -4460 4238 -4356 4362
rect -4460 4222 -4333 4238
rect -8489 4110 -4567 4111
rect -8489 190 -8488 4110
rect -4568 190 -4567 4110
rect -8489 189 -4567 190
rect -6580 -189 -6476 189
rect -4460 78 -4413 4222
rect -4349 78 -4333 4222
rect -2261 4111 -2157 4489
rect -141 4378 -94 8522
rect -30 4378 -14 8522
rect 2058 8411 2162 8600
rect 4178 8538 4282 8600
rect 4178 8522 4305 8538
rect 149 8410 4071 8411
rect 149 4490 150 8410
rect 4070 4490 4071 8410
rect 149 4489 4071 4490
rect -141 4362 -14 4378
rect -141 4238 -37 4362
rect -141 4222 -14 4238
rect -4170 4110 -248 4111
rect -4170 190 -4169 4110
rect -249 190 -248 4110
rect -4170 189 -248 190
rect -4460 62 -4333 78
rect -4460 -62 -4356 62
rect -4460 -78 -4333 -62
rect -8489 -190 -4567 -189
rect -8489 -4110 -8488 -190
rect -4568 -4110 -4567 -190
rect -8489 -4111 -4567 -4110
rect -6580 -4489 -6476 -4111
rect -4460 -4222 -4413 -78
rect -4349 -4222 -4333 -78
rect -2261 -189 -2157 189
rect -141 78 -94 4222
rect -30 78 -14 4222
rect 2058 4111 2162 4489
rect 4178 4378 4225 8522
rect 4289 4378 4305 8522
rect 6377 8411 6481 8600
rect 8497 8538 8601 8600
rect 8497 8522 8624 8538
rect 4468 8410 8390 8411
rect 4468 4490 4469 8410
rect 8389 4490 8390 8410
rect 4468 4489 8390 4490
rect 4178 4362 4305 4378
rect 4178 4238 4282 4362
rect 4178 4222 4305 4238
rect 149 4110 4071 4111
rect 149 190 150 4110
rect 4070 190 4071 4110
rect 149 189 4071 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -4170 -190 -248 -189
rect -4170 -4110 -4169 -190
rect -249 -4110 -248 -190
rect -4170 -4111 -248 -4110
rect -4460 -4238 -4333 -4222
rect -4460 -4362 -4356 -4238
rect -4460 -4378 -4333 -4362
rect -8489 -4490 -4567 -4489
rect -8489 -8410 -8488 -4490
rect -4568 -8410 -4567 -4490
rect -8489 -8411 -4567 -8410
rect -6580 -8600 -6476 -8411
rect -4460 -8522 -4413 -4378
rect -4349 -8522 -4333 -4378
rect -2261 -4489 -2157 -4111
rect -141 -4222 -94 -78
rect -30 -4222 -14 -78
rect 2058 -189 2162 189
rect 4178 78 4225 4222
rect 4289 78 4305 4222
rect 6377 4111 6481 4489
rect 8497 4378 8544 8522
rect 8608 4378 8624 8522
rect 8497 4362 8624 4378
rect 8497 4238 8601 4362
rect 8497 4222 8624 4238
rect 4468 4110 8390 4111
rect 4468 190 4469 4110
rect 8389 190 8390 4110
rect 4468 189 8390 190
rect 4178 62 4305 78
rect 4178 -62 4282 62
rect 4178 -78 4305 -62
rect 149 -190 4071 -189
rect 149 -4110 150 -190
rect 4070 -4110 4071 -190
rect 149 -4111 4071 -4110
rect -141 -4238 -14 -4222
rect -141 -4362 -37 -4238
rect -141 -4378 -14 -4362
rect -4170 -4490 -248 -4489
rect -4170 -8410 -4169 -4490
rect -249 -8410 -248 -4490
rect -4170 -8411 -248 -8410
rect -4460 -8538 -4333 -8522
rect -4460 -8600 -4356 -8538
rect -2261 -8600 -2157 -8411
rect -141 -8522 -94 -4378
rect -30 -8522 -14 -4378
rect 2058 -4489 2162 -4111
rect 4178 -4222 4225 -78
rect 4289 -4222 4305 -78
rect 6377 -189 6481 189
rect 8497 78 8544 4222
rect 8608 78 8624 4222
rect 8497 62 8624 78
rect 8497 -62 8601 62
rect 8497 -78 8624 -62
rect 4468 -190 8390 -189
rect 4468 -4110 4469 -190
rect 8389 -4110 8390 -190
rect 4468 -4111 8390 -4110
rect 4178 -4238 4305 -4222
rect 4178 -4362 4282 -4238
rect 4178 -4378 4305 -4362
rect 149 -4490 4071 -4489
rect 149 -8410 150 -4490
rect 4070 -8410 4071 -4490
rect 149 -8411 4071 -8410
rect -141 -8538 -14 -8522
rect -141 -8600 -37 -8538
rect 2058 -8600 2162 -8411
rect 4178 -8522 4225 -4378
rect 4289 -8522 4305 -4378
rect 6377 -4489 6481 -4111
rect 8497 -4222 8544 -78
rect 8608 -4222 8624 -78
rect 8497 -4238 8624 -4222
rect 8497 -4362 8601 -4238
rect 8497 -4378 8624 -4362
rect 4468 -4490 8390 -4489
rect 4468 -8410 4469 -4490
rect 8389 -8410 8390 -4490
rect 4468 -8411 8390 -8410
rect 4178 -8538 4305 -8522
rect 4178 -8600 4282 -8538
rect 6377 -8600 6481 -8411
rect 8497 -8522 8544 -4378
rect 8608 -8522 8624 -4378
rect 8497 -8538 8624 -8522
rect 8497 -8600 8601 -8538
<< properties >>
string FIXED_BBOX 4329 4350 8529 8550
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 20 l 20 val 815.2 carea 2.00 cperi 0.19 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
