magic
tech sky130A
magscale 1 2
timestamp 1725111581
<< viali >>
rect 11092 -4506 19992 -4472
rect 11092 -5014 19426 -4980
rect 11092 -5106 19426 -5072
rect 11690 -5614 19992 -5580
rect 11690 -5706 19992 -5672
<< metal1 >>
rect 1590 6620 2270 10320
rect 1590 4980 2280 5680
rect 1590 1170 2260 1870
rect 1590 -600 2260 800
rect 20250 -910 20700 -900
rect 20250 -1560 20260 -910
rect 20690 -1560 20700 -910
rect 10960 -4340 11550 -4110
rect 15530 -4340 15770 -4130
rect 19560 -4340 20160 -4140
rect 10960 -4472 20160 -4340
rect 10960 -4506 11092 -4472
rect 19992 -4506 20160 -4472
rect 10960 -4520 20160 -4506
rect 10960 -4970 11550 -4520
rect 10960 -4980 19454 -4970
rect 10960 -5014 11092 -4980
rect 19426 -5014 19454 -4980
rect 1590 -5650 10670 -5020
rect 10250 -5820 10670 -5650
rect 10960 -5072 19454 -5014
rect 10960 -5106 11092 -5072
rect 19426 -5106 19454 -5072
rect 10960 -5120 19454 -5106
rect 10960 -5710 11080 -5120
rect 11140 -5820 11550 -5210
rect 19531 -5474 19952 -4611
rect 20045 -5570 20160 -4520
rect 11640 -5580 20160 -5570
rect 11640 -5614 11690 -5580
rect 19992 -5614 20160 -5580
rect 11640 -5672 20160 -5614
rect 11640 -5706 11690 -5672
rect 19992 -5706 20160 -5672
rect 11640 -5710 20160 -5706
rect 11640 -5720 20070 -5710
rect 20250 -5820 20700 -1560
rect 10250 -6070 11550 -5820
rect 19570 -6070 20700 -5820
rect 20250 -6380 20700 -6070
rect 19430 -7020 20700 -6380
<< via1 >>
rect 20260 -1560 20690 -910
<< metal2 >>
rect 1590 -4740 2870 -3880
use ldoota  ldoota_0
timestamp 1724262930
transform 1 0 3650 0 1 1170
box -1490 -8480 17521 9150
use sky130_fd_pr__res_xhigh_po_1p41_4KNYXQ  sky130_fd_pr__res_xhigh_po_1p41_4KNYXQ_0
timestamp 1725111581
transform 0 1 15542 -1 0 -4743
box -307 -4582 307 4582
use sky130_fd_pr__res_xhigh_po_1p41_4KNYXQ  sky130_fd_pr__res_xhigh_po_1p41_4KNYXQ_1
timestamp 1725111581
transform 0 1 15542 -1 0 -5943
box -307 -4582 307 4582
use sky130_fd_pr__res_xhigh_po_1p41_4KNYXQ  sky130_fd_pr__res_xhigh_po_1p41_4KNYXQ_2
timestamp 1725111581
transform 0 1 15542 -1 0 -5343
box -307 -4582 307 4582
<< labels >>
flabel metal1 19430 -7020 20700 -6380 0 FreeSans 1600 0 0 0 VLDO
port 4 nsew
flabel metal1 1590 -5650 2060 -5020 0 FreeSans 1600 0 0 0 FBOUT
port 6 nsew
flabel metal1 1590 1170 2060 1870 0 FreeSans 1600 0 0 0 FBIN
port 5 nsew
flabel metal1 1590 -600 2060 800 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal2 1590 -4740 2060 -3880 0 FreeSans 1600 0 0 0 IB
port 2 nsew
flabel metal1 1590 4980 2060 5680 0 FreeSans 1600 0 0 0 VREF
port 3 nsew
flabel metal1 1590 6620 2060 10320 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
<< end >>
