magic
tech sky130A
magscale 1 2
timestamp 1725202727
<< nwell >>
rect 3413 3230 4051 3264
rect 181 880 861 1134
rect 452 735 486 769
rect 3867 568 4174 1134
<< pwell >>
rect 3457 2414 4174 2799
rect -1004 2014 -352 2048
rect -306 1536 3380 1550
rect 3439 1536 4174 2414
rect -306 1332 4174 1536
rect -299 259 3830 334
<< psubdiff >>
rect 4067 2508 4134 2539
rect -1004 2014 -352 2048
rect 4067 1577 4074 2508
rect 4128 1577 4134 2508
rect 4067 1542 4134 1577
rect -310 296 3830 299
rect -310 262 -274 296
rect 3791 262 3830 296
rect -310 259 3830 262
<< nsubdiff >>
rect 3413 3230 4051 3264
rect 330 1002 617 1032
rect 330 900 362 1002
rect 578 900 617 1002
rect 330 869 617 900
rect 3865 863 4138 868
rect 3865 808 3894 863
rect 4095 808 4138 863
rect 3865 803 4138 808
<< psubdiffcont >>
rect 4074 1577 4128 2508
rect -274 262 3791 296
<< nsubdiffcont >>
rect 362 900 578 1002
rect 3894 808 4095 863
<< locali >>
rect 4067 2508 4135 2539
rect 4067 1577 4074 2508
rect 4128 1577 4135 2508
rect 4067 1541 4135 1577
rect 330 1002 617 1032
rect 330 900 362 1002
rect 578 900 617 1002
rect 330 834 617 900
rect 3828 863 4174 868
rect 3828 808 3894 863
rect 4095 808 4174 863
rect 3828 803 4174 808
rect -310 296 3830 324
rect -310 262 -274 296
rect 3791 262 3830 296
rect -310 259 3830 262
<< viali >>
rect -279 3230 4051 3264
rect -1004 2014 -352 2048
rect -270 1572 3310 1606
rect 4074 1577 4128 2508
rect -284 1060 -240 1169
rect -187 1136 118 1174
rect 914 1146 965 1251
rect 1034 1145 1325 1179
rect 1364 1146 1432 1180
rect 1742 1130 1817 1196
rect 1926 1146 1960 1180
rect 2012 1146 2046 1180
rect 3742 1078 3812 1200
rect 362 915 578 1002
rect 3494 936 3559 970
rect 421 735 486 769
rect 1921 664 1972 766
rect 2261 732 2326 766
rect 3761 664 3812 766
rect -281 529 -8 563
rect 80 452 114 622
rect 168 502 238 624
rect 2008 502 2078 624
<< metal1 >>
rect -315 3346 4147 3361
rect -315 3228 -298 3346
rect 377 3264 4147 3346
rect 4051 3230 4147 3264
rect 377 3228 4147 3230
rect -315 3212 4147 3228
rect -58 3110 266 3212
rect 674 3110 998 3212
rect 1406 3110 1730 3212
rect 2138 3110 2462 3212
rect 2870 3110 3194 3212
rect 3602 3110 3926 3212
rect -183 3082 -96 3100
rect 304 3082 636 3100
rect 1036 3082 1368 3100
rect 1768 3082 2100 3100
rect 2500 3082 2832 3100
rect 3232 3082 3564 3100
rect 3964 3082 4051 3100
rect -183 3026 4051 3082
rect -183 3008 -96 3026
rect 304 3008 636 3026
rect 1036 3008 1368 3026
rect 1768 3008 2100 3026
rect 2500 3008 2832 3026
rect 3232 3008 4051 3026
rect -888 2982 -367 2998
rect -888 2847 -490 2982
rect -383 2847 -367 2982
rect -888 2832 -367 2847
rect -888 2666 -564 2832
rect -58 2724 266 2998
rect 674 2724 998 2998
rect 1406 2724 1730 2998
rect 2138 2724 2462 2998
rect 2870 2724 3194 2998
rect 3477 2952 4051 3008
rect -183 2696 -96 2714
rect 304 2696 391 2714
rect -1216 2638 -926 2656
rect -526 2638 -448 2656
rect -1216 2582 -448 2638
rect -183 2640 391 2696
rect -183 2622 -96 2640
rect 304 2622 391 2640
rect 549 2696 636 2714
rect 1036 2696 1123 2714
rect 549 2640 1123 2696
rect 549 2622 636 2640
rect 1036 2622 1123 2640
rect 1281 2696 1368 2714
rect 1768 2696 1855 2714
rect 1281 2640 1855 2696
rect 1281 2622 1368 2640
rect 1768 2622 1855 2640
rect 2013 2696 2100 2714
rect 2500 2696 2587 2714
rect 2013 2640 2587 2696
rect 2013 2622 2100 2640
rect 2500 2622 2587 2640
rect 2745 2696 2832 2714
rect 3232 2696 3319 2714
rect 2745 2640 3319 2696
rect 3602 2686 3926 2952
rect 2745 2622 2832 2640
rect 3232 2622 3319 2640
rect 3460 2658 3564 2676
rect 3964 2658 4183 2812
rect -1216 2564 -926 2582
rect -526 2564 -448 2582
rect -1216 1254 -1157 2564
rect -888 2458 -564 2554
rect -174 2458 -128 2622
rect -888 2378 -128 2458
rect -888 2280 -564 2378
rect -1126 2252 -926 2270
rect -526 2252 -448 2270
rect -1126 2196 -448 2252
rect -1126 2178 -926 2196
rect -526 2178 -448 2196
rect -174 2214 -128 2378
rect -58 2458 266 2612
rect 558 2458 604 2622
rect -58 2378 604 2458
rect -58 2224 266 2378
rect 558 2214 604 2378
rect 674 2458 998 2612
rect 1290 2458 1336 2622
rect 674 2378 1336 2458
rect 674 2224 998 2378
rect 1290 2214 1336 2378
rect 1406 2458 1730 2612
rect 2022 2458 2068 2622
rect 1406 2449 2068 2458
rect 1406 2387 1415 2449
rect 1721 2387 2068 2449
rect 1406 2378 2068 2387
rect 1406 2224 1730 2378
rect 2022 2214 2068 2378
rect 2138 2458 2462 2612
rect 2754 2458 2800 2622
rect 2138 2378 2800 2458
rect 2138 2224 2462 2378
rect 2754 2214 2800 2378
rect 2870 2451 3194 2612
rect 2870 2384 2877 2451
rect 3187 2384 3194 2451
rect 2870 2224 3194 2384
rect 3460 2602 4183 2658
rect 3460 2584 3564 2602
rect 3964 2585 4183 2602
rect 3964 2584 4042 2585
rect 3460 2295 3532 2584
rect 3602 2553 3926 2574
rect 3602 2508 4175 2553
rect 3602 2407 4074 2508
rect 3460 2249 3664 2295
rect -174 2196 -96 2214
rect 304 2196 382 2214
rect -1126 1348 -1063 2178
rect -888 2060 -564 2168
rect -174 2140 382 2196
rect -174 2122 -96 2140
rect 304 2122 382 2140
rect 558 2196 636 2214
rect 1036 2196 1114 2214
rect 558 2140 1114 2196
rect 558 2122 636 2140
rect 1036 2122 1114 2140
rect 1290 2196 1368 2214
rect 1768 2196 1846 2214
rect 1290 2140 1846 2196
rect 1290 2122 1368 2140
rect 1768 2122 1846 2140
rect 2022 2196 2100 2214
rect 2500 2196 2578 2214
rect 2022 2140 2578 2196
rect 2022 2122 2100 2140
rect 2500 2122 2578 2140
rect 2754 2196 2832 2214
rect 3232 2196 3310 2214
rect 2754 2140 3310 2196
rect 2754 2122 2832 2140
rect 3232 2122 3310 2140
rect -1015 2048 -226 2060
rect -1015 2014 -1004 2048
rect -352 2014 -226 2048
rect -1015 1962 -226 2014
rect -1015 1806 -999 1962
rect -703 1806 -226 1962
rect -58 1838 266 2112
rect 674 1838 998 2112
rect 1406 1838 1730 2112
rect 2138 1838 2462 2112
rect 2870 1838 3194 2112
rect 3460 1979 3617 2249
rect 3963 2137 4074 2407
rect 3867 2091 4074 2137
rect 3460 1933 3665 1979
rect 3460 1828 3617 1933
rect -1015 1791 -226 1806
rect -352 1627 -226 1791
rect -174 1810 -96 1828
rect 304 1810 636 1828
rect 1036 1810 1368 1828
rect 1768 1810 2100 1828
rect 2500 1810 2832 1828
rect 3232 1810 3617 1828
rect 3963 1821 4074 2091
rect -174 1754 3617 1810
rect 3858 1775 4074 1821
rect -174 1736 -96 1754
rect 304 1736 636 1754
rect 1036 1736 1368 1754
rect 1768 1736 2100 1754
rect 2500 1736 2832 1754
rect 3232 1736 3617 1754
rect -58 1627 266 1726
rect 674 1627 998 1726
rect 1406 1627 1730 1726
rect 2138 1627 2462 1726
rect 2870 1627 3194 1726
rect 3263 1673 3617 1736
rect 3460 1663 3617 1673
rect -352 1606 3380 1627
rect 3460 1617 3667 1663
rect -352 1572 -270 1606
rect 3310 1577 3380 1606
rect 3963 1577 4074 1775
rect 4128 1577 4175 2508
rect 3310 1572 4175 1577
rect -352 1519 4175 1572
rect -1126 1314 -404 1348
rect -352 1347 4174 1519
rect -1126 1285 983 1314
rect -1216 1217 863 1254
rect -1216 1191 -379 1217
rect -316 1169 -231 1186
rect -316 1128 -284 1169
rect -1218 1060 -284 1128
rect -240 1060 -231 1169
rect -203 1174 138 1180
rect -203 1166 -187 1174
rect 118 1166 138 1174
rect -203 1094 -189 1166
rect 123 1094 138 1166
rect -203 1081 138 1094
rect 178 1135 777 1182
rect -1218 1053 -231 1060
rect 178 1053 219 1135
rect 650 1102 694 1103
rect -1218 999 219 1053
rect 255 1062 694 1102
rect 255 967 299 1062
rect -429 927 299 967
rect 330 1002 617 1032
rect -429 775 -348 927
rect 330 915 362 1002
rect 578 915 617 1002
rect 650 967 694 1062
rect 731 1031 777 1135
rect 813 1104 863 1217
rect 897 1251 983 1285
rect 897 1146 914 1251
rect 965 1146 983 1251
rect 1577 1266 2181 1309
rect 897 1139 983 1146
rect 1015 1196 1319 1197
rect 1015 1180 1441 1196
rect 1015 1179 1364 1180
rect 1015 1145 1034 1179
rect 1325 1146 1364 1179
rect 1432 1146 1441 1180
rect 1325 1145 1441 1146
rect 1015 1130 1441 1145
rect 1015 1104 1340 1130
rect 813 1066 1340 1104
rect 1577 1099 1679 1266
rect 1374 1031 1679 1099
rect 731 999 1679 1031
rect 1730 1196 1829 1202
rect 1730 1130 1742 1196
rect 1817 1130 1829 1196
rect 1917 1180 2053 1196
rect 1917 1146 1926 1180
rect 1960 1146 2012 1180
rect 2046 1146 2053 1180
rect 1917 1130 2053 1146
rect 1730 1007 1829 1130
rect 2097 1102 2181 1266
rect 2301 1235 4033 1304
rect 3730 1200 3830 1206
rect 3730 1102 3742 1200
rect 2097 1078 3742 1102
rect 3812 1102 3830 1200
rect 3812 1078 3970 1102
rect 2097 1072 3970 1078
rect 1730 967 1830 1007
rect 650 927 1830 967
rect 3482 970 3571 976
rect 3482 936 3494 970
rect 3559 967 3571 970
rect 3559 936 3904 967
rect 3482 930 3904 936
rect 330 891 617 915
rect -1215 769 498 775
rect 3865 772 3904 930
rect -1215 735 421 769
rect 486 735 498 769
rect -1215 734 498 735
rect -1215 681 143 734
rect 409 729 498 734
rect 1909 766 2338 772
rect 1909 664 1921 766
rect 1972 735 2261 766
rect 1972 664 1984 735
rect 2249 732 2261 735
rect 2326 732 2338 766
rect 2249 726 2338 732
rect 3749 766 3904 772
rect 1909 658 1984 664
rect 3749 664 3761 766
rect 3812 664 3904 766
rect 3749 658 3904 664
rect 68 622 126 644
rect 3940 630 3970 1072
rect -1216 575 -314 602
rect -1216 563 6 575
rect -1216 529 -281 563
rect -8 529 6 563
rect -1216 517 6 529
rect -1216 481 -314 517
rect 68 452 80 622
rect 114 467 126 622
rect 156 624 3970 630
rect 156 502 168 624
rect 238 600 2008 624
rect 238 502 250 600
rect 156 496 250 502
rect 1990 502 2008 600
rect 2078 600 3970 624
rect 2078 502 2090 600
rect 1990 496 2090 502
rect 4000 467 4033 1235
rect 114 452 4033 467
rect 68 398 4033 452
rect 4069 355 4174 1347
rect 3820 259 4174 355
<< via1 >>
rect -298 3264 377 3346
rect -298 3230 -279 3264
rect -279 3230 377 3264
rect -298 3228 377 3230
rect -490 2847 -383 2982
rect 1415 2387 1721 2449
rect 2877 2384 3187 2451
rect -999 1806 -703 1962
rect -189 1136 -187 1166
rect -187 1136 118 1166
rect 118 1136 123 1166
rect -189 1094 123 1136
rect -300 813 141 889
<< metal2 >>
rect -1216 3361 -506 3362
rect -1216 3346 392 3361
rect -1216 3228 -298 3346
rect 377 3228 392 3346
rect -1216 3212 392 3228
rect -1216 1962 -690 1974
rect -1216 1806 -999 1962
rect -703 1806 -690 1962
rect -1216 1791 -690 1806
rect -662 899 -535 3212
rect -506 2982 3194 2998
rect -506 2847 -490 2982
rect -383 2847 3194 2982
rect -506 2832 3194 2847
rect 1406 2449 1730 2458
rect 1406 2387 1415 2449
rect 1721 2387 1730 2449
rect 1406 1180 1730 2387
rect 2870 2451 3194 2832
rect 2870 2384 2877 2451
rect 3187 2384 3194 2451
rect 2870 2378 3194 2384
rect -202 1166 1730 1180
rect -202 1094 -189 1166
rect 123 1094 1730 1166
rect -202 1081 1730 1094
rect -662 889 227 899
rect -662 813 -300 889
rect 141 813 227 889
rect -662 803 227 813
use sky130_fd_pr__nfet_01v8_AXXKZX  sky130_fd_pr__nfet_01v8_AXXKZX_0
timestamp 1642872912
transform 0 1 104 -1 0 2168
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_AXXKZX  sky130_fd_pr__nfet_01v8_AXXKZX_1
timestamp 1642872912
transform 0 1 104 -1 0 1782
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_AXXKZX  sky130_fd_pr__nfet_01v8_AXXKZX_2
timestamp 1642872912
transform 0 1 836 -1 0 2168
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_AXXKZX  sky130_fd_pr__nfet_01v8_AXXKZX_3
timestamp 1642872912
transform 0 1 836 -1 0 1782
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_AXXKZX  sky130_fd_pr__nfet_01v8_AXXKZX_4
timestamp 1642872912
transform 0 1 3032 -1 0 1782
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_AXXKZX  sky130_fd_pr__nfet_01v8_AXXKZX_5
timestamp 1642872912
transform 0 1 2300 -1 0 1782
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_AXXKZX  sky130_fd_pr__nfet_01v8_AXXKZX_6
timestamp 1642872912
transform 0 1 2300 -1 0 2168
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_AXXKZX  sky130_fd_pr__nfet_01v8_AXXKZX_7
timestamp 1642872912
transform 0 1 3032 -1 0 2168
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_AXXKZX  sky130_fd_pr__nfet_01v8_AXXKZX_8
timestamp 1642872912
transform 0 1 1568 -1 0 1782
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_AXXKZX  sky130_fd_pr__nfet_01v8_AXXKZX_9
timestamp 1642872912
transform 0 1 1568 -1 0 2168
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_AXXKZX  sky130_fd_pr__nfet_01v8_AXXKZX_10
timestamp 1642872912
transform 0 1 -726 -1 0 2224
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_AXXKZX  sky130_fd_pr__nfet_01v8_AXXKZX_11
timestamp 1642872912
transform 0 1 -726 -1 0 2610
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_HS2QBX  sky130_fd_pr__nfet_01v8_HS2QBX_0
timestamp 1642973952
transform 0 1 3764 -1 0 2630
box -108 -288 108 288
use sky130_fd_pr__nfet_01v8_HW54L5  sky130_fd_pr__nfet_01v8_HW54L5_0
timestamp 1642973952
transform 0 1 3733 -1 0 2035
box -424 -257 424 257
use sky130_fd_pr__pfet_01v8_9ZL4AL  sky130_fd_pr__pfet_01v8_9ZL4AL_0
timestamp 1642872912
transform 0 1 104 -1 0 2668
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_9ZL4AL  sky130_fd_pr__pfet_01v8_9ZL4AL_1
timestamp 1642872912
transform 0 1 104 -1 0 3054
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_9ZL4AL  sky130_fd_pr__pfet_01v8_9ZL4AL_2
timestamp 1642872912
transform 0 1 836 -1 0 3054
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_9ZL4AL  sky130_fd_pr__pfet_01v8_9ZL4AL_3
timestamp 1642872912
transform 0 1 836 -1 0 2668
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_9ZL4AL  sky130_fd_pr__pfet_01v8_9ZL4AL_4
timestamp 1642872912
transform 0 1 2300 -1 0 3054
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_9ZL4AL  sky130_fd_pr__pfet_01v8_9ZL4AL_5
timestamp 1642872912
transform 0 1 2300 -1 0 2668
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_9ZL4AL  sky130_fd_pr__pfet_01v8_9ZL4AL_6
timestamp 1642872912
transform 0 1 3032 -1 0 2668
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_9ZL4AL  sky130_fd_pr__pfet_01v8_9ZL4AL_7
timestamp 1642872912
transform 0 1 1568 -1 0 2668
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_9ZL4AL  sky130_fd_pr__pfet_01v8_9ZL4AL_8
timestamp 1642872912
transform 0 1 1568 -1 0 3054
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_9ZL4AL  sky130_fd_pr__pfet_01v8_9ZL4AL_9
timestamp 1642872912
transform 0 1 3032 -1 0 3054
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_9ZL4AL  sky130_fd_pr__pfet_01v8_9ZL4AL_10
timestamp 1642872912
transform 0 1 3764 -1 0 3054
box -246 -419 246 419
use sky130_fd_sc_hd__dfrtn_1  sky130_fd_sc_hd__dfrtn_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 150 0 1 307
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtn_1  sky130_fd_sc_hd__dfrtn_1_1
timestamp 1723858470
transform 1 0 1990 0 1 307
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtn_1  sky130_fd_sc_hd__dfrtn_1_3
timestamp 1723858470
transform -1 0 3830 0 -1 1395
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 -310 0 1 307
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_1
timestamp 1723858470
transform -1 0 150 0 -1 1395
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_2
timestamp 1723858470
transform -1 0 1346 0 -1 1395
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  sky130_fd_sc_hd__or2_4_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 1990 0 -1 1395
box -38 -48 682 592
<< labels >>
flabel metal2 -1216 1791 -1126 1974 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel metal1 -1218 999 -1123 1128 0 FreeSans 800 0 0 0 OSC
port 6 nsew
flabel metal1 -1215 681 -1120 775 0 FreeSans 800 0 0 0 EN
port 4 nsew
flabel metal1 -1216 481 -1121 602 0 FreeSans 800 0 0 0 RESET
port 5 nsew
flabel metal2 -1216 3213 -1124 3362 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel metal1 3713 948 3713 948 0 FreeSans 320 0 0 0 ENA_D1
flabel metal1 4094 2585 4183 2812 0 FreeSans 1600 0 0 0 IB
port 3 nsew
<< end >>
