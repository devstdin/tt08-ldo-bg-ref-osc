magic
tech sky130A
magscale 1 2
timestamp 1725107840
<< nwell >>
rect -950 1150 3600 1840
rect -950 -6500 5030 1150
<< pwell >>
rect -1820 3280 9170 3660
rect -1820 -6500 -950 3280
rect 3600 1150 9170 3280
rect 5030 -6500 9170 1150
rect -1820 -9510 9170 -6500
<< mvpsubdiff >>
rect -1180 -6640 5220 -6620
rect -1180 -6710 70 -6640
rect 4070 -6710 5220 -6640
rect -1180 -6730 5220 -6710
rect -1180 -6830 -1070 -6730
rect -1180 -8790 -1160 -6830
rect -1090 -8790 -1070 -6830
rect -1180 -8870 -1070 -8790
rect 5110 -6830 5220 -6730
rect 5110 -8790 5130 -6830
rect 5200 -8790 5220 -6830
rect 5110 -8870 5220 -8790
rect -1180 -8890 5220 -8870
rect -1180 -8960 70 -8890
rect 4070 -8960 5220 -8890
rect -1180 -8980 5220 -8960
<< mvnsubdiff >>
rect -850 1030 4930 1050
rect -850 970 70 1030
rect 4070 970 4930 1030
rect -850 950 4930 970
rect -850 770 -750 950
rect -850 -6140 -830 770
rect -770 -6140 -750 770
rect -850 -6300 -750 -6140
rect 4830 770 4930 950
rect 4830 -6140 4850 770
rect 4910 -6140 4930 770
rect 4830 -6300 4930 -6140
rect -850 -6320 4930 -6300
rect -850 -6380 70 -6320
rect 4070 -6380 4930 -6320
rect -850 -6400 4930 -6380
<< mvpsubdiffcont >>
rect 70 -6710 4070 -6640
rect -1160 -8790 -1090 -6830
rect 5130 -8790 5200 -6830
rect 70 -8960 4070 -8890
<< mvnsubdiffcont >>
rect 70 970 4070 1030
rect -830 -6140 -770 770
rect 4850 -6140 4910 770
rect 70 -6380 4070 -6320
<< locali >>
rect -830 970 70 1030
rect 4070 970 4910 1030
rect -830 770 -770 970
rect -830 -6320 -770 -6140
rect 4850 770 4910 970
rect 4850 -6320 4910 -6140
rect -830 -6380 70 -6320
rect 4070 -6380 4910 -6320
rect -1160 -6710 70 -6640
rect 4070 -6710 5200 -6640
rect -1160 -6830 -1090 -6710
rect -1160 -8890 -1090 -8790
rect 5130 -6830 5200 -6710
rect 5130 -8890 5200 -8790
rect -1160 -8960 70 -8890
rect 4070 -8960 5200 -8890
<< viali >>
rect -776 3162 -208 3196
rect -50 3162 518 3196
rect 676 3162 1244 3196
rect 1402 3162 1970 3196
rect 2128 3162 2696 3196
rect 2854 3162 3422 3196
rect -776 1758 -208 1792
rect 70 970 4070 1030
rect -830 -6140 -770 770
rect 4850 -6140 4910 770
rect 7554 -6268 7588 -5918
rect 70 -6380 4070 -6320
rect 5192 -6364 7492 -6330
rect 70 -6710 4070 -6640
rect -1160 -8790 -1090 -6830
rect 5130 -8790 5200 -6830
rect 70 -8960 4070 -8890
rect 8672 -8936 8706 -7708
rect 5474 -9032 6042 -8998
rect 6330 -9032 6898 -8998
rect 7186 -9032 7754 -8998
rect 8042 -9032 8610 -8998
<< metal1 >>
rect -1820 3650 3600 3660
rect -1820 3160 -1660 3650
rect -990 3196 3600 3650
rect -990 3162 -776 3196
rect -208 3162 -50 3196
rect 518 3162 676 3196
rect 1244 3162 1402 3196
rect 1970 3162 2128 3196
rect 2696 3162 2854 3196
rect 3422 3162 3600 3196
rect -990 3160 3600 3162
rect -1820 3150 3600 3160
rect -790 3020 -290 3100
rect -790 2880 -720 3020
rect -1820 2370 -700 2880
rect -1670 2250 -980 2260
rect -1670 1790 -1660 2250
rect -990 1800 -980 2250
rect -790 2070 -700 2370
rect -590 2660 -390 3020
rect -260 2980 -180 3150
rect -590 2360 -580 2660
rect -400 2360 -390 2660
rect -790 1940 -720 2070
rect -590 1940 -390 2360
rect -290 2070 -180 2980
rect -70 2980 0 3150
rect -70 2070 20 2980
rect 140 2660 340 3050
rect 140 2360 150 2660
rect 330 2360 340 2660
rect -790 1858 -290 1940
rect 140 1900 340 2360
rect 440 2070 750 2880
rect 860 2660 1060 3050
rect 1190 2980 1260 3150
rect 860 2360 870 2660
rect 1050 2360 1060 2660
rect -990 1792 -100 1800
rect -990 1790 -776 1792
rect -1670 1758 -776 1790
rect -208 1758 -100 1792
rect -1670 1040 -100 1758
rect 490 1310 700 2070
rect 860 1900 1060 2360
rect 1170 2070 1260 2980
rect 1390 2980 1460 3150
rect 1390 2070 1480 2980
rect 1590 2660 1790 3050
rect 2110 2980 2180 3150
rect 1590 2360 1600 2660
rect 1780 2360 1790 2660
rect 1590 1900 1790 2360
rect 1890 1980 2070 2880
rect 2110 2070 2200 2980
rect 2310 2660 2510 3050
rect 2840 2980 2910 3150
rect 2310 2360 2320 2660
rect 2500 2360 2510 2660
rect 1910 1840 2070 1980
rect 2310 1900 2510 2360
rect 2620 1980 2790 2880
rect 2840 2070 2930 2980
rect 3040 2660 3240 3050
rect 3040 2360 3050 2660
rect 3230 2360 3240 2660
rect 2640 1840 2790 1980
rect 3040 1900 3240 2360
rect 3350 2690 3520 2880
rect 3350 2050 9170 2690
rect 1910 1820 2790 1840
rect 3390 1820 9170 2050
rect 1910 1440 9170 1820
rect 490 1110 500 1310
rect 690 1110 700 1310
rect 490 1100 700 1110
rect 5130 1160 8330 1170
rect -1670 1030 4920 1040
rect -1670 970 70 1030
rect 4070 970 4920 1030
rect -1670 770 4920 970
rect -1670 -6140 -830 770
rect -770 460 4850 770
rect -770 -5830 -630 460
rect -546 348 4402 400
rect 4524 348 4695 400
rect 70 329 4070 348
rect -547 166 -538 283
rect -425 166 4695 283
rect -17 165 4157 166
rect 70 100 4070 118
rect -546 99 4070 100
rect -546 47 4226 99
rect 4348 47 4695 99
rect -546 14 4695 15
rect -546 -38 -385 14
rect -263 -37 4695 14
rect -263 -38 4070 -37
rect 70 -56 4070 -38
rect -17 -106 4157 -105
rect -546 -223 4573 -106
rect 4689 -223 4695 -106
rect 70 -288 4070 -270
rect -546 -289 4070 -288
rect -546 -341 -219 -289
rect -97 -341 4695 -289
rect -546 -427 4226 -375
rect 4348 -427 4695 -375
rect -546 -428 4070 -427
rect 70 -446 4070 -428
rect -17 -494 4157 -493
rect -547 -611 -538 -494
rect -425 -611 4695 -494
rect 70 -676 4070 -658
rect -546 -677 4070 -676
rect -546 -729 4402 -677
rect 4524 -729 4695 -677
rect -546 -764 4695 -763
rect -546 -816 -219 -764
rect -97 -815 4695 -764
rect -97 -816 4070 -815
rect 70 -834 4070 -816
rect -17 -882 4157 -881
rect -546 -999 4573 -882
rect 4689 -999 4695 -882
rect 70 -1064 4070 -1046
rect -546 -1065 4070 -1064
rect -546 -1117 -385 -1065
rect -263 -1117 4695 -1065
rect -546 -1203 4402 -1151
rect 4524 -1203 4695 -1151
rect -546 -1204 4070 -1203
rect 70 -1222 4070 -1204
rect -17 -1270 4157 -1269
rect -547 -1387 -538 -1270
rect -425 -1387 4695 -1270
rect 70 -1452 4070 -1434
rect -546 -1453 4070 -1452
rect -546 -1505 4226 -1453
rect 4348 -1505 4695 -1453
rect -546 -1540 4695 -1539
rect -546 -1592 -385 -1540
rect -263 -1591 4695 -1540
rect -263 -1592 4070 -1591
rect 70 -1610 4070 -1592
rect -17 -1658 4157 -1657
rect -546 -1775 4573 -1658
rect 4689 -1775 4695 -1658
rect 70 -1840 4070 -1822
rect -546 -1841 4070 -1840
rect -546 -1893 -219 -1841
rect -97 -1893 4695 -1841
rect -546 -1979 4226 -1927
rect 4348 -1979 4695 -1927
rect -546 -1980 4070 -1979
rect 70 -1998 4070 -1980
rect -17 -2046 4157 -2045
rect -547 -2163 -538 -2046
rect -425 -2163 4695 -2046
rect 70 -2228 4070 -2210
rect -546 -2229 4070 -2228
rect -546 -2281 4402 -2229
rect 4524 -2281 4695 -2229
rect -546 -2316 4695 -2315
rect -546 -2368 -219 -2316
rect -97 -2367 4695 -2316
rect -97 -2368 4070 -2367
rect 70 -2386 4070 -2368
rect -17 -2434 4157 -2433
rect -546 -2551 4573 -2434
rect 4689 -2551 4695 -2434
rect 70 -2616 4070 -2598
rect -546 -2617 4070 -2616
rect -546 -2669 -385 -2617
rect -263 -2669 4695 -2617
rect -546 -2704 4695 -2703
rect -546 -2756 -385 -2704
rect -263 -2755 4695 -2704
rect -263 -2756 4070 -2755
rect 70 -2774 4070 -2756
rect -17 -2822 4157 -2821
rect -546 -2939 4573 -2822
rect 4689 -2939 4695 -2822
rect 70 -3004 4070 -2986
rect -546 -3005 4070 -3004
rect -546 -3057 -219 -3005
rect -97 -3057 4695 -3005
rect -546 -3143 4402 -3091
rect 4524 -3143 4695 -3091
rect -546 -3144 4070 -3143
rect 70 -3162 4070 -3144
rect -17 -3210 4157 -3209
rect -547 -3327 -538 -3210
rect -425 -3327 4695 -3210
rect 70 -3392 4070 -3374
rect -546 -3393 4070 -3392
rect -546 -3445 4226 -3393
rect 4348 -3445 4695 -3393
rect -546 -3480 4695 -3479
rect -546 -3532 -219 -3480
rect -97 -3531 4695 -3480
rect -97 -3532 4070 -3531
rect 70 -3550 4070 -3532
rect -17 -3598 4157 -3597
rect -546 -3715 4573 -3598
rect 4689 -3715 4695 -3598
rect 70 -3780 4070 -3762
rect -546 -3781 4070 -3780
rect -546 -3833 -385 -3781
rect -263 -3833 4695 -3781
rect -546 -3919 4226 -3867
rect 4348 -3919 4695 -3867
rect -546 -3920 4070 -3919
rect 70 -3938 4070 -3920
rect -17 -3986 4157 -3985
rect -547 -4103 -538 -3986
rect -425 -4103 4695 -3986
rect 70 -4168 4070 -4150
rect -546 -4169 4070 -4168
rect -546 -4221 4402 -4169
rect 4524 -4221 4695 -4169
rect -546 -4256 4695 -4255
rect -546 -4308 -385 -4256
rect -263 -4307 4695 -4256
rect -263 -4308 4070 -4307
rect 70 -4326 4070 -4308
rect -17 -4374 4157 -4373
rect -546 -4491 4573 -4374
rect 4689 -4491 4695 -4374
rect 70 -4556 4070 -4538
rect -546 -4557 4070 -4556
rect -546 -4609 -219 -4557
rect -97 -4609 4695 -4557
rect -546 -4695 4402 -4643
rect 4524 -4695 4695 -4643
rect -546 -4696 4070 -4695
rect 70 -4714 4070 -4696
rect -17 -4762 4157 -4761
rect -547 -4879 -538 -4762
rect -425 -4879 4695 -4762
rect 70 -4944 4070 -4926
rect -546 -4945 4070 -4944
rect -546 -4997 4226 -4945
rect 4348 -4997 4695 -4945
rect -546 -5032 4695 -5031
rect -546 -5084 -219 -5032
rect -97 -5083 4695 -5032
rect -97 -5084 4070 -5083
rect 70 -5102 4070 -5084
rect -17 -5150 4157 -5149
rect -546 -5267 4573 -5150
rect 4689 -5267 4695 -5150
rect 70 -5332 4070 -5314
rect -546 -5333 4070 -5332
rect -546 -5385 -385 -5333
rect -263 -5385 4695 -5333
rect -546 -5471 4226 -5419
rect 4348 -5471 4695 -5419
rect -546 -5472 4070 -5471
rect 70 -5490 4070 -5472
rect -17 -5538 4157 -5537
rect -547 -5655 -538 -5538
rect -425 -5655 4695 -5538
rect 70 -5720 4070 -5702
rect -546 -5721 4070 -5720
rect -546 -5773 4402 -5721
rect 4524 -5773 4695 -5721
rect 4750 -5830 4850 460
rect -770 -6140 4850 -5830
rect 4910 -6140 4920 770
rect 5130 700 5140 1160
rect 8320 700 8330 1160
rect 5130 690 8330 700
rect 6530 -5754 7500 690
rect -1670 -6320 4920 -6140
rect 5150 -5850 5760 -5830
rect 5150 -6260 5170 -5850
rect 5730 -6260 5760 -5850
rect 6530 -6240 7468 -5754
rect 7543 -5918 7700 -5897
rect 5150 -6280 5760 -6260
rect 7543 -6268 7554 -5918
rect 7588 -6268 7700 -5918
rect 7543 -6320 7700 -6268
rect -1670 -6380 70 -6320
rect 4070 -6380 4920 -6320
rect -1670 -6390 4920 -6380
rect 4990 -6330 7700 -6320
rect 4990 -6364 5192 -6330
rect 7492 -6364 7700 -6330
rect 4990 -6500 7700 -6364
rect -1670 -6640 5330 -6500
rect -1670 -6710 70 -6640
rect 4070 -6710 5330 -6640
rect -1670 -6740 5330 -6710
rect -1670 -6830 -320 -6740
rect 1350 -6830 1400 -6740
rect 2630 -6830 2680 -6740
rect 4350 -6830 5330 -6740
rect -1670 -8790 -1160 -6830
rect -1090 -6960 -320 -6830
rect -210 -6840 50 -6830
rect -210 -6920 -200 -6840
rect 40 -6920 50 -6840
rect -1090 -6970 -270 -6960
rect -1090 -7050 -360 -6970
rect -280 -7050 -270 -6970
rect -1090 -7060 -270 -7050
rect -1090 -7190 -320 -7060
rect -1090 -8430 -435 -7190
rect -370 -7246 -334 -7190
rect -370 -7310 -320 -7246
rect -370 -8310 -300 -7310
rect -370 -8374 -320 -8310
rect -370 -8430 -334 -8374
rect -1090 -8440 -320 -8430
rect -1090 -8520 -540 -8440
rect -330 -8520 -320 -8440
rect -1090 -8790 -320 -8520
rect -210 -8700 50 -6920
rect 150 -7090 200 -6830
rect 100 -7100 200 -7090
rect 100 -7180 110 -7100
rect 190 -7180 200 -7100
rect 100 -7190 200 -7180
rect 150 -7310 200 -7190
rect 130 -8310 200 -7310
rect -210 -8780 -200 -8700
rect 40 -8780 50 -8700
rect -210 -8790 50 -8780
rect 150 -8790 200 -8310
rect 230 -6840 330 -6830
rect 230 -6920 240 -6840
rect 320 -6920 330 -6840
rect 230 -6930 330 -6920
rect 390 -6840 650 -6830
rect 390 -6920 400 -6840
rect 640 -6920 650 -6840
rect 230 -7310 280 -6930
rect 230 -8310 310 -7310
rect 230 -8560 280 -8310
rect 230 -8570 330 -8560
rect 230 -8650 240 -8570
rect 320 -8650 330 -8570
rect 230 -8660 330 -8650
rect 390 -8570 650 -6920
rect 750 -7310 800 -6830
rect 730 -8310 800 -7310
rect 750 -8430 800 -8310
rect 700 -8440 800 -8430
rect 700 -8520 710 -8440
rect 790 -8520 800 -8440
rect 700 -8530 800 -8520
rect 390 -8650 400 -8570
rect 640 -8650 650 -8570
rect 230 -8690 280 -8660
rect 230 -8700 330 -8690
rect 230 -8780 240 -8700
rect 320 -8780 330 -8700
rect 230 -8790 330 -8780
rect 390 -8700 650 -8650
rect 390 -8780 400 -8700
rect 640 -8780 650 -8700
rect 390 -8790 650 -8780
rect -1670 -8850 -320 -8790
rect 750 -8850 800 -8530
rect 830 -7090 880 -6830
rect 990 -6840 1250 -6830
rect 990 -6920 1000 -6840
rect 1240 -6920 1250 -6840
rect 830 -7100 930 -7090
rect 830 -7180 840 -7100
rect 920 -7180 930 -7100
rect 830 -7190 930 -7180
rect 830 -7310 880 -7190
rect 830 -8310 910 -7310
rect 830 -8790 880 -8310
rect 990 -8700 1250 -6920
rect 1350 -6960 1480 -6830
rect 1300 -6970 1480 -6960
rect 1300 -7050 1310 -6970
rect 1390 -7050 1480 -6970
rect 1300 -7060 1480 -7050
rect 1350 -7310 1480 -7060
rect 1580 -6840 1840 -6830
rect 1580 -6920 1590 -6840
rect 1830 -6920 1840 -6840
rect 1330 -8310 1510 -7310
rect 990 -8780 1000 -8700
rect 1240 -8780 1250 -8700
rect 990 -8790 1250 -8780
rect 1350 -8430 1480 -8310
rect 1350 -8440 1530 -8430
rect 1350 -8520 1440 -8440
rect 1520 -8520 1530 -8440
rect 1350 -8530 1530 -8520
rect 1350 -8850 1480 -8530
rect 1580 -8570 1840 -6920
rect 1900 -6840 2000 -6830
rect 1900 -6920 1910 -6840
rect 1990 -6920 2000 -6840
rect 1900 -6930 2000 -6920
rect 1950 -7310 2000 -6930
rect 1930 -8310 2000 -7310
rect 1950 -8560 2000 -8310
rect 1580 -8650 1590 -8570
rect 1830 -8650 1840 -8570
rect 1580 -8700 1840 -8650
rect 1900 -8570 2000 -8560
rect 1900 -8650 1910 -8570
rect 1990 -8650 2000 -8570
rect 1900 -8660 2000 -8650
rect 1950 -8690 2000 -8660
rect 1580 -8780 1590 -8700
rect 1830 -8780 1840 -8700
rect 1580 -8790 1840 -8780
rect 1900 -8700 2000 -8690
rect 1900 -8780 1910 -8700
rect 1990 -8780 2000 -8700
rect 1900 -8790 2000 -8780
rect 2030 -6840 2130 -6830
rect 2030 -6920 2040 -6840
rect 2120 -6920 2130 -6840
rect 2030 -6930 2130 -6920
rect 2190 -6840 2450 -6830
rect 2190 -6920 2200 -6840
rect 2440 -6920 2450 -6840
rect 2030 -7310 2080 -6930
rect 2030 -8310 2100 -7310
rect 2030 -8560 2080 -8310
rect 2030 -8570 2130 -8560
rect 2030 -8650 2040 -8570
rect 2120 -8650 2130 -8570
rect 2030 -8660 2130 -8650
rect 2190 -8570 2450 -6920
rect 2550 -6960 2680 -6830
rect 2790 -6840 3050 -6830
rect 2790 -6920 2800 -6840
rect 3040 -6920 3050 -6840
rect 2550 -6970 2730 -6960
rect 2550 -7050 2640 -6970
rect 2720 -7050 2730 -6970
rect 2550 -7060 2730 -7050
rect 2550 -7310 2680 -7060
rect 2530 -8310 2700 -7310
rect 2550 -8430 2680 -8310
rect 2500 -8440 2680 -8430
rect 2500 -8520 2510 -8440
rect 2590 -8520 2680 -8440
rect 2500 -8530 2680 -8520
rect 2190 -8650 2200 -8570
rect 2440 -8650 2450 -8570
rect 2030 -8690 2080 -8660
rect 2030 -8700 2130 -8690
rect 2030 -8780 2040 -8700
rect 2120 -8780 2130 -8700
rect 2030 -8790 2130 -8780
rect 2190 -8700 2450 -8650
rect 2190 -8780 2200 -8700
rect 2440 -8780 2450 -8700
rect 2190 -8790 2450 -8780
rect 2550 -8850 2680 -8530
rect 2790 -8700 3050 -6920
rect 3150 -7090 3200 -6830
rect 3100 -7100 3200 -7090
rect 3100 -7180 3110 -7100
rect 3190 -7180 3200 -7100
rect 3100 -7190 3200 -7180
rect 3150 -7310 3200 -7190
rect 3130 -8310 3200 -7310
rect 2790 -8780 2800 -8700
rect 3040 -8780 3050 -8700
rect 2790 -8790 3050 -8780
rect 3150 -8790 3200 -8310
rect 3230 -7310 3280 -6830
rect 3380 -6840 3640 -6830
rect 3380 -6920 3390 -6840
rect 3630 -6920 3640 -6840
rect 3230 -8310 3310 -7310
rect 3230 -8430 3280 -8310
rect 3230 -8440 3330 -8430
rect 3230 -8520 3240 -8440
rect 3320 -8520 3330 -8440
rect 3230 -8530 3330 -8520
rect 3230 -8850 3280 -8530
rect 3380 -8570 3640 -6920
rect 3700 -6840 3800 -6830
rect 3700 -6920 3710 -6840
rect 3790 -6920 3800 -6840
rect 3700 -6930 3800 -6920
rect 3750 -7310 3800 -6930
rect 3730 -8310 3800 -7310
rect 3750 -8560 3800 -8310
rect 3380 -8650 3390 -8570
rect 3630 -8650 3640 -8570
rect 3380 -8700 3640 -8650
rect 3700 -8570 3800 -8560
rect 3700 -8650 3710 -8570
rect 3790 -8650 3800 -8570
rect 3700 -8660 3800 -8650
rect 3750 -8690 3800 -8660
rect 3380 -8780 3390 -8700
rect 3630 -8780 3640 -8700
rect 3380 -8790 3640 -8780
rect 3700 -8700 3800 -8690
rect 3700 -8780 3710 -8700
rect 3790 -8780 3800 -8700
rect 3700 -8790 3800 -8780
rect 3830 -7090 3880 -6830
rect 3990 -6840 4250 -6830
rect 3990 -6920 4000 -6840
rect 4240 -6920 4250 -6840
rect 3830 -7100 3930 -7090
rect 3830 -7180 3840 -7100
rect 3920 -7180 3930 -7100
rect 3830 -7190 3930 -7180
rect 3830 -7310 3880 -7190
rect 3830 -8310 3910 -7310
rect 3830 -8790 3880 -8310
rect 3990 -8700 4250 -6920
rect 4350 -6960 5130 -6830
rect 4300 -6970 5130 -6960
rect 4300 -7050 4310 -6970
rect 4390 -7050 5130 -6970
rect 4300 -7060 5130 -7050
rect 4330 -8312 4404 -7310
rect 4343 -8425 4404 -8312
rect 4460 -8425 5130 -7060
rect 4343 -8440 5130 -8425
rect 4343 -8520 4375 -8440
rect 4560 -8520 5130 -8440
rect 4343 -8530 5130 -8520
rect 3990 -8780 4000 -8700
rect 4240 -8780 4250 -8700
rect 3990 -8790 4250 -8780
rect 4370 -8790 5130 -8530
rect 5200 -7690 5330 -6830
rect 5460 -6540 5550 -6530
rect 5460 -6830 5470 -6540
rect 5540 -6830 5550 -6540
rect 5200 -8790 5400 -7690
rect 5460 -7710 5550 -6830
rect 5650 -6890 5870 -6530
rect 5650 -7180 5660 -6890
rect 5860 -7180 5870 -6890
rect 5460 -7820 5530 -7710
rect 5460 -8730 5550 -7820
rect 4370 -8850 5400 -8790
rect -1820 -8890 5400 -8850
rect -1820 -8960 70 -8890
rect 4070 -8960 5400 -8890
rect 5650 -8900 5870 -7180
rect 5970 -7240 6060 -6530
rect 5970 -7530 5980 -7240
rect 6050 -7530 6060 -7240
rect 5970 -7710 6060 -7530
rect 5990 -7820 6060 -7710
rect 5970 -8730 6060 -7820
rect 6310 -6540 6400 -6530
rect 6310 -6830 6320 -6540
rect 6390 -6830 6400 -6540
rect 6310 -7710 6400 -6830
rect 6510 -6890 6730 -6530
rect 6510 -7180 6520 -6890
rect 6720 -7180 6730 -6890
rect 6310 -7820 6380 -7710
rect 6310 -8730 6400 -7820
rect 6510 -8900 6730 -7180
rect 6820 -7240 6910 -6530
rect 6820 -7530 6830 -7240
rect 6900 -7530 6910 -7240
rect 6820 -7710 6910 -7530
rect 6840 -7820 6910 -7710
rect 6820 -8730 6910 -7820
rect 7170 -6540 7260 -6530
rect 7170 -6830 7180 -6540
rect 7250 -6830 7260 -6540
rect 7170 -7710 7260 -6830
rect 7360 -6890 7580 -6530
rect 7360 -7180 7370 -6890
rect 7570 -7180 7580 -6890
rect 7170 -7820 7240 -7710
rect 7170 -8730 7260 -7820
rect 7360 -8900 7580 -7180
rect 7680 -7240 7770 -6530
rect 7680 -7530 7690 -7240
rect 7760 -7530 7770 -7240
rect 7680 -7710 7770 -7530
rect 7700 -7820 7770 -7710
rect 7680 -8730 7770 -7820
rect 8030 -6540 8120 -6530
rect 8030 -6830 8040 -6540
rect 8110 -6830 8120 -6540
rect 8030 -7710 8120 -6830
rect 8210 -6890 8430 -6530
rect 8580 -6540 9170 1440
rect 8580 -6830 8590 -6540
rect 9160 -6830 9170 -6540
rect 8580 -6850 9170 -6830
rect 8210 -7180 8220 -6890
rect 8420 -7180 8430 -6890
rect 8030 -7820 8100 -7710
rect 8030 -8730 8120 -7820
rect 8210 -8900 8430 -7180
rect 8540 -7240 9170 -7230
rect 8540 -7530 8550 -7240
rect 8620 -7530 9170 -7240
rect 8540 -7540 9170 -7530
rect 8540 -7710 8630 -7540
rect 8670 -7702 9170 -7540
rect 8560 -7820 8630 -7710
rect 8540 -8730 8630 -7820
rect 8665 -7708 9170 -7702
rect 8665 -8936 8672 -7708
rect 8706 -8936 9170 -7708
rect 8665 -8947 9170 -8936
rect -1820 -8980 5400 -8960
rect 8670 -8980 9170 -8947
rect -1820 -8998 9170 -8980
rect -1820 -9032 5474 -8998
rect 6042 -9032 6330 -8998
rect 6898 -9032 7186 -8998
rect 7754 -9032 8042 -8998
rect 8610 -9032 9170 -8998
rect -1820 -9510 9170 -9032
<< via1 >>
rect -1660 3160 -990 3650
rect -1660 1790 -990 2250
rect -580 2360 -400 2660
rect 150 2360 330 2660
rect 870 2360 1050 2660
rect 1600 2360 1780 2660
rect 2320 2360 2500 2660
rect 3050 2360 3230 2660
rect 500 1110 690 1310
rect 4402 348 4524 400
rect -538 166 -425 283
rect 4226 47 4348 99
rect -385 -38 -263 14
rect 4573 -223 4689 -106
rect -219 -341 -97 -289
rect 4226 -427 4348 -375
rect -538 -611 -425 -494
rect 4402 -729 4524 -677
rect -219 -816 -97 -764
rect 4573 -999 4689 -882
rect -385 -1117 -263 -1065
rect 4402 -1203 4524 -1151
rect -538 -1387 -425 -1270
rect 4226 -1505 4348 -1453
rect -385 -1592 -263 -1540
rect 4573 -1775 4689 -1658
rect -219 -1893 -97 -1841
rect 4226 -1979 4348 -1927
rect -538 -2163 -425 -2046
rect 4402 -2281 4524 -2229
rect -219 -2368 -97 -2316
rect 4573 -2551 4689 -2434
rect -385 -2669 -263 -2617
rect -385 -2756 -263 -2704
rect 4573 -2939 4689 -2822
rect -219 -3057 -97 -3005
rect 4402 -3143 4524 -3091
rect -538 -3327 -425 -3210
rect 4226 -3445 4348 -3393
rect -219 -3532 -97 -3480
rect 4573 -3715 4689 -3598
rect -385 -3833 -263 -3781
rect 4226 -3919 4348 -3867
rect -538 -4103 -425 -3986
rect 4402 -4221 4524 -4169
rect -385 -4308 -263 -4256
rect 4573 -4491 4689 -4374
rect -219 -4609 -97 -4557
rect 4402 -4695 4524 -4643
rect -538 -4879 -425 -4762
rect 4226 -4997 4348 -4945
rect -219 -5084 -97 -5032
rect 4573 -5267 4689 -5150
rect -385 -5385 -263 -5333
rect 4226 -5471 4348 -5419
rect -538 -5655 -425 -5538
rect 4402 -5773 4524 -5721
rect 5140 700 8320 1160
rect 5170 -6260 5730 -5850
rect -200 -6920 40 -6840
rect -360 -7050 -280 -6970
rect -540 -8520 -330 -8440
rect 110 -7180 190 -7100
rect -200 -8780 40 -8700
rect 240 -6920 320 -6840
rect 400 -6920 640 -6840
rect 240 -8650 320 -8570
rect 710 -8520 790 -8440
rect 400 -8650 640 -8570
rect 240 -8780 320 -8700
rect 400 -8780 640 -8700
rect 1000 -6920 1240 -6840
rect 840 -7180 920 -7100
rect 1310 -7050 1390 -6970
rect 1590 -6920 1830 -6840
rect 1000 -8780 1240 -8700
rect 1440 -8520 1520 -8440
rect 1910 -6920 1990 -6840
rect 1590 -8650 1830 -8570
rect 1910 -8650 1990 -8570
rect 1590 -8780 1830 -8700
rect 1910 -8780 1990 -8700
rect 2040 -6920 2120 -6840
rect 2200 -6920 2440 -6840
rect 2040 -8650 2120 -8570
rect 2800 -6920 3040 -6840
rect 2640 -7050 2720 -6970
rect 2510 -8520 2590 -8440
rect 2200 -8650 2440 -8570
rect 2040 -8780 2120 -8700
rect 2200 -8780 2440 -8700
rect 3110 -7180 3190 -7100
rect 2800 -8780 3040 -8700
rect 3390 -6920 3630 -6840
rect 3240 -8520 3320 -8440
rect 3710 -6920 3790 -6840
rect 3390 -8650 3630 -8570
rect 3710 -8650 3790 -8570
rect 3390 -8780 3630 -8700
rect 3710 -8780 3790 -8700
rect 4000 -6920 4240 -6840
rect 3840 -7180 3920 -7100
rect 4310 -7050 4390 -6970
rect 4375 -8520 4560 -8440
rect 4000 -8780 4240 -8700
rect 5470 -6830 5540 -6540
rect 5660 -7180 5860 -6890
rect 5980 -7530 6050 -7240
rect 6320 -6830 6390 -6540
rect 6520 -7180 6720 -6890
rect 6830 -7530 6900 -7240
rect 7180 -6830 7250 -6540
rect 7370 -7180 7570 -6890
rect 7690 -7530 7760 -7240
rect 8040 -6830 8110 -6540
rect 8590 -6830 9160 -6540
rect 8220 -7180 8420 -6890
rect 8550 -7530 8620 -7240
<< metal2 >>
rect -1670 3650 -980 3660
rect -1670 3160 -1660 3650
rect -990 3160 -980 3650
rect -1670 2250 -980 3160
rect -590 2660 3250 2670
rect -590 2360 -580 2660
rect -400 2360 150 2660
rect 330 2360 870 2660
rect 1050 2360 1600 2660
rect 1780 2360 2320 2660
rect 2500 2360 3050 2660
rect 3230 2360 3250 2660
rect -590 2350 3250 2360
rect -1670 1790 -1660 2250
rect -990 1790 -980 2250
rect -1670 1780 -980 1790
rect -1820 1390 1790 1650
rect -1820 1130 360 1390
rect 820 1320 1790 1390
rect 490 1310 700 1320
rect 490 1110 500 1310
rect 690 1110 700 1310
rect 820 1130 4700 1320
rect 490 1060 700 1110
rect -220 810 4350 1060
rect -550 283 -420 300
rect -550 166 -538 283
rect -425 166 -420 283
rect -550 50 -420 166
rect -1820 -490 -420 50
rect -550 -494 -420 -490
rect -550 -611 -538 -494
rect -425 -611 -420 -494
rect -550 -1270 -420 -611
rect -550 -1387 -538 -1270
rect -425 -1387 -420 -1270
rect -550 -2046 -420 -1387
rect -550 -2163 -538 -2046
rect -425 -2163 -420 -2046
rect -550 -3210 -420 -2163
rect -550 -3327 -538 -3210
rect -425 -3327 -420 -3210
rect -550 -3986 -420 -3327
rect -550 -4103 -538 -3986
rect -425 -4103 -420 -3986
rect -550 -4762 -420 -4103
rect -550 -4879 -538 -4762
rect -425 -4879 -420 -4762
rect -550 -5538 -420 -4879
rect -550 -5655 -538 -5538
rect -425 -5655 -420 -5538
rect -550 -5670 -420 -5655
rect -390 14 -260 30
rect -390 -38 -385 14
rect -263 -38 -260 14
rect -390 -1065 -260 -38
rect -390 -1117 -385 -1065
rect -263 -1117 -260 -1065
rect -390 -1540 -260 -1117
rect -390 -1592 -385 -1540
rect -263 -1592 -260 -1540
rect -390 -2617 -260 -1592
rect -390 -2669 -385 -2617
rect -263 -2669 -260 -2617
rect -390 -2704 -260 -2669
rect -390 -2756 -385 -2704
rect -263 -2756 -260 -2704
rect -390 -3781 -260 -2756
rect -390 -3833 -385 -3781
rect -263 -3833 -260 -3781
rect -390 -4256 -260 -3833
rect -390 -4308 -385 -4256
rect -263 -4308 -260 -4256
rect -390 -5333 -260 -4308
rect -220 -289 -90 810
rect -220 -341 -219 -289
rect -97 -341 -90 -289
rect -220 -764 -90 -341
rect -220 -816 -219 -764
rect -97 -816 -90 -764
rect -220 -1841 -90 -816
rect -220 -1893 -219 -1841
rect -97 -1893 -90 -1841
rect -220 -2316 -90 -1893
rect -220 -2368 -219 -2316
rect -97 -2368 -90 -2316
rect -220 -3005 -90 -2368
rect -220 -3057 -219 -3005
rect -97 -3057 -90 -3005
rect -220 -3480 -90 -3057
rect -220 -3532 -219 -3480
rect -97 -3532 -90 -3480
rect -220 -4557 -90 -3532
rect -220 -4609 -219 -4557
rect -97 -4609 -90 -4557
rect -220 -5032 -90 -4609
rect -220 -5084 -219 -5032
rect -97 -5084 -90 -5032
rect -220 -5100 -90 -5084
rect 4220 99 4350 810
rect 4400 470 4700 1130
rect 5130 1160 8330 1170
rect 5130 700 5140 1160
rect 8320 700 8330 1160
rect 5130 690 8330 700
rect 4220 47 4226 99
rect 4348 47 4350 99
rect 4220 -375 4350 47
rect 4220 -427 4226 -375
rect 4348 -427 4350 -375
rect 4220 -1453 4350 -427
rect 4220 -1505 4226 -1453
rect 4348 -1505 4350 -1453
rect 4220 -1927 4350 -1505
rect 4220 -1979 4226 -1927
rect 4348 -1979 4350 -1927
rect 4220 -3393 4350 -1979
rect 4220 -3445 4226 -3393
rect 4348 -3445 4350 -3393
rect 4220 -3867 4350 -3445
rect 4220 -3919 4226 -3867
rect 4348 -3919 4350 -3867
rect 4220 -4945 4350 -3919
rect 4220 -4997 4226 -4945
rect 4348 -4997 4350 -4945
rect -390 -5385 -385 -5333
rect -263 -5385 -260 -5333
rect -390 -5720 -260 -5385
rect 4220 -5419 4350 -4997
rect 4220 -5471 4226 -5419
rect 4348 -5471 4350 -5419
rect 4220 -5490 4350 -5471
rect 4400 400 4530 410
rect 4400 348 4402 400
rect 4524 348 4530 400
rect 4400 -677 4530 348
rect 4400 -729 4402 -677
rect 4524 -729 4530 -677
rect 4400 -1151 4530 -729
rect 4400 -1203 4402 -1151
rect 4524 -1203 4530 -1151
rect 4400 -2229 4530 -1203
rect 4400 -2281 4402 -2229
rect 4524 -2281 4530 -2229
rect 4400 -3091 4530 -2281
rect 4400 -3143 4402 -3091
rect 4524 -3143 4530 -3091
rect 4400 -4169 4530 -3143
rect 4400 -4221 4402 -4169
rect 4524 -4221 4530 -4169
rect 4400 -4643 4530 -4221
rect 4400 -4695 4402 -4643
rect 4524 -4695 4530 -4643
rect 4400 -5490 4530 -4695
rect 4570 -106 4700 470
rect 4570 -223 4573 -106
rect 4689 -223 4700 -106
rect 4570 -882 4700 -223
rect 4570 -999 4573 -882
rect 4689 -999 4700 -882
rect 4570 -1658 4700 -999
rect 4570 -1775 4573 -1658
rect 4689 -1775 4700 -1658
rect 4570 -2434 4700 -1775
rect 4570 -2551 4573 -2434
rect 4689 -2551 4700 -2434
rect 4570 -2822 4700 -2551
rect 4570 -2939 4573 -2822
rect 4689 -2939 4700 -2822
rect 4570 -3598 4700 -2939
rect 4570 -3715 4573 -3598
rect 4689 -3715 4700 -3598
rect 4570 -4374 4700 -3715
rect 4570 -4491 4573 -4374
rect 4689 -4491 4700 -4374
rect 4570 -5150 4700 -4491
rect 4570 -5267 4573 -5150
rect 4689 -5267 4700 -5150
rect 4570 -5290 4700 -5267
rect -550 -6770 -90 -5720
rect 4400 -5721 4800 -5490
rect 4400 -5773 4402 -5721
rect 4524 -5773 4800 -5721
rect 4400 -5830 4800 -5773
rect 4400 -5850 5760 -5830
rect 4400 -6260 5170 -5850
rect 5730 -6260 5760 -5850
rect 4400 -6280 5760 -6260
rect 7770 -5920 8330 -5900
rect 4400 -6360 4940 -6280
rect 4400 -6700 4800 -6360
rect 7770 -6380 7790 -5920
rect 8310 -6380 8330 -5920
rect 7770 -6530 8330 -6380
rect -550 -6840 4430 -6770
rect -550 -6920 -200 -6840
rect 40 -6920 240 -6840
rect 320 -6920 400 -6840
rect 640 -6920 1000 -6840
rect 1240 -6920 1590 -6840
rect 1830 -6920 1910 -6840
rect 1990 -6920 2040 -6840
rect 2120 -6920 2200 -6840
rect 2440 -6920 2800 -6840
rect 3040 -6920 3390 -6840
rect 3630 -6920 3710 -6840
rect 3790 -6920 4000 -6840
rect 4240 -6920 4430 -6840
rect -550 -6930 4430 -6920
rect 4500 -6880 4800 -6700
rect 5400 -6540 9170 -6530
rect 5400 -6830 5470 -6540
rect 5540 -6830 6320 -6540
rect 6390 -6830 7180 -6540
rect 7250 -6830 8040 -6540
rect 8110 -6830 8590 -6540
rect 9160 -6830 9170 -6540
rect 5400 -6840 9170 -6830
rect 4500 -6890 8430 -6880
rect -400 -6970 4430 -6960
rect -400 -7050 -360 -6970
rect -280 -7050 1310 -6970
rect 1390 -7050 2640 -6970
rect 2720 -7050 4310 -6970
rect 4390 -7050 4430 -6970
rect -400 -7060 4430 -7050
rect 4500 -7090 5660 -6890
rect -400 -7100 5660 -7090
rect -400 -7180 110 -7100
rect 190 -7180 840 -7100
rect 920 -7180 3110 -7100
rect 3190 -7180 3840 -7100
rect 3920 -7180 5660 -7100
rect 5860 -7180 6520 -6890
rect 6720 -7180 7370 -6890
rect 7570 -7180 8220 -6890
rect 8420 -7180 8430 -6890
rect -400 -7190 8430 -7180
rect 5400 -7240 8630 -7230
rect 5400 -7530 5980 -7240
rect 6050 -7530 6830 -7240
rect 6900 -7530 7690 -7240
rect 7760 -7530 8550 -7240
rect 8620 -7530 8630 -7240
rect 5400 -7540 8630 -7530
rect -550 -8440 4570 -8430
rect -550 -8520 -540 -8440
rect -330 -8520 710 -8440
rect 790 -8520 1440 -8440
rect 1520 -8520 2510 -8440
rect 2590 -8520 3240 -8440
rect 3320 -8520 4375 -8440
rect 4560 -8520 4570 -8440
rect -550 -8530 4570 -8520
rect -400 -8570 4430 -8560
rect -400 -8650 240 -8570
rect 320 -8650 400 -8570
rect 640 -8650 1590 -8570
rect 1830 -8650 1910 -8570
rect 1990 -8650 2040 -8570
rect 2120 -8650 2200 -8570
rect 2440 -8650 3390 -8570
rect 3630 -8650 3710 -8570
rect 3790 -8650 4430 -8570
rect -400 -8660 4430 -8650
rect -400 -8700 4430 -8690
rect -400 -8780 -200 -8700
rect 40 -8780 240 -8700
rect 320 -8780 400 -8700
rect 640 -8780 1000 -8700
rect 1240 -8780 1590 -8700
rect 1830 -8780 1910 -8700
rect 1990 -8780 2040 -8700
rect 2120 -8780 2200 -8700
rect 2440 -8780 2800 -8700
rect 3040 -8780 3390 -8700
rect 3630 -8780 3710 -8700
rect 3790 -8780 4000 -8700
rect 4240 -8780 4430 -8700
rect -400 -8790 4430 -8780
<< via2 >>
rect 5170 730 8290 1130
rect 7790 -6380 8310 -5920
<< metal3 >>
rect 5130 1130 8330 1170
rect 5130 730 5170 1130
rect 8290 730 8330 1130
rect 5130 690 8330 730
rect 7770 -5920 8330 -5460
rect 7770 -6380 7790 -5920
rect 8310 -6380 8330 -5920
rect 7770 -6400 8330 -6380
<< via3 >>
rect 5220 780 8240 1080
<< metal4 >>
rect 5130 1080 8330 1170
rect 5130 780 5220 1080
rect 8240 780 8330 1080
rect 5130 -5620 8330 780
use sky130_fd_pr__cap_mim_m3_1_5WMUWD  sky130_fd_pr__cap_mim_m3_1_5WMUWD_0
timestamp 1646668631
transform 1 0 6780 0 1 -2620
box -1750 -3100 1749 3100
use sky130_fd_pr__nfet_g5v0d10v5_DP5JSB  sky130_fd_pr__nfet_g5v0d10v5_DP5JSB_0
timestamp 1646652369
transform 1 0 -682 0 1 -7812
box -258 -588 258 588
use sky130_fd_pr__nfet_g5v0d10v5_DP5JSB  sky130_fd_pr__nfet_g5v0d10v5_DP5JSB_1
timestamp 1646652369
transform 1 0 -82 0 1 -7812
box -258 -588 258 588
use sky130_fd_pr__nfet_g5v0d10v5_DP5JSB  sky130_fd_pr__nfet_g5v0d10v5_DP5JSB_2
timestamp 1646652369
transform 1 0 518 0 1 -7812
box -258 -588 258 588
use sky130_fd_pr__nfet_g5v0d10v5_DP5JSB  sky130_fd_pr__nfet_g5v0d10v5_DP5JSB_3
timestamp 1646652369
transform 1 0 1118 0 1 -7812
box -258 -588 258 588
use sky130_fd_pr__nfet_g5v0d10v5_DP5JSB  sky130_fd_pr__nfet_g5v0d10v5_DP5JSB_4
timestamp 1646652369
transform 1 0 1718 0 1 -7812
box -258 -588 258 588
use sky130_fd_pr__nfet_g5v0d10v5_DP5JSB  sky130_fd_pr__nfet_g5v0d10v5_DP5JSB_5
timestamp 1646652369
transform 1 0 2318 0 1 -7812
box -258 -588 258 588
use sky130_fd_pr__nfet_g5v0d10v5_DP5JSB  sky130_fd_pr__nfet_g5v0d10v5_DP5JSB_6
timestamp 1646652369
transform 1 0 2918 0 1 -7812
box -258 -588 258 588
use sky130_fd_pr__nfet_g5v0d10v5_DP5JSB  sky130_fd_pr__nfet_g5v0d10v5_DP5JSB_7
timestamp 1646652369
transform 1 0 3518 0 1 -7812
box -258 -588 258 588
use sky130_fd_pr__nfet_g5v0d10v5_DP5JSB  sky130_fd_pr__nfet_g5v0d10v5_DP5JSB_8
timestamp 1646652369
transform 1 0 4118 0 1 -7812
box -258 -588 258 588
use sky130_fd_pr__nfet_g5v0d10v5_DP5JSB  sky130_fd_pr__nfet_g5v0d10v5_DP5JSB_9
timestamp 1646652369
transform 1 0 4718 0 1 -7812
box -258 -588 258 588
use sky130_fd_pr__nfet_g5v0d10v5_RQRC42  sky130_fd_pr__nfet_g5v0d10v5_RQRC42_0
timestamp 1646668631
transform 1 0 5758 0 1 -8322
box -428 -758 428 758
use sky130_fd_pr__nfet_g5v0d10v5_RQRC42  sky130_fd_pr__nfet_g5v0d10v5_RQRC42_1
timestamp 1646668631
transform 1 0 6614 0 1 -8322
box -428 -758 428 758
use sky130_fd_pr__nfet_g5v0d10v5_RQRC42  sky130_fd_pr__nfet_g5v0d10v5_RQRC42_2
timestamp 1646668631
transform 1 0 7470 0 1 -8322
box -428 -758 428 758
use sky130_fd_pr__nfet_g5v0d10v5_RQRC42  sky130_fd_pr__nfet_g5v0d10v5_RQRC42_3
timestamp 1646668631
transform 1 0 8326 0 1 -8322
box -428 -758 428 758
use sky130_fd_pr__pfet_g5v0d10v5_JNK3YL  sky130_fd_pr__pfet_g5v0d10v5_JNK3YL_0
timestamp 1646668020
transform 1 0 -492 0 1 2477
box -458 -797 458 797
use sky130_fd_pr__pfet_g5v0d10v5_JNK3YL  sky130_fd_pr__pfet_g5v0d10v5_JNK3YL_1
timestamp 1646668020
transform 1 0 234 0 1 2477
box -458 -797 458 797
use sky130_fd_pr__pfet_g5v0d10v5_JNK3YL  sky130_fd_pr__pfet_g5v0d10v5_JNK3YL_2
timestamp 1646668020
transform 1 0 960 0 1 2477
box -458 -797 458 797
use sky130_fd_pr__pfet_g5v0d10v5_JNK3YL  sky130_fd_pr__pfet_g5v0d10v5_JNK3YL_3
timestamp 1646668020
transform 1 0 1686 0 1 2477
box -458 -797 458 797
use sky130_fd_pr__pfet_g5v0d10v5_JNK3YL  sky130_fd_pr__pfet_g5v0d10v5_JNK3YL_4
timestamp 1646668020
transform 1 0 2412 0 1 2477
box -458 -797 458 797
use sky130_fd_pr__pfet_g5v0d10v5_JNK3YL  sky130_fd_pr__pfet_g5v0d10v5_JNK3YL_5
timestamp 1646668020
transform 1 0 3138 0 1 2477
box -458 -797 458 797
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_0
timestamp 1646595912
transform 0 1 2070 -1 0 224
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_1
timestamp 1646595912
transform 0 1 2070 -1 0 -164
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_2
timestamp 1646595912
transform 0 1 2070 -1 0 -552
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_3
timestamp 1646595912
transform 0 1 2070 -1 0 -940
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_4
timestamp 1646595912
transform 0 1 2070 -1 0 -1328
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_5
timestamp 1646595912
transform 0 1 2070 -1 0 -1716
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_6
timestamp 1646595912
transform 0 1 2070 -1 0 -2104
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_7
timestamp 1646595912
transform 0 1 2070 -1 0 -2492
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_8
timestamp 1646595912
transform 0 1 2070 -1 0 -2880
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_9
timestamp 1646595912
transform 0 1 2070 -1 0 -3268
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_10
timestamp 1646595912
transform 0 1 2070 -1 0 -3656
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_11
timestamp 1646595912
transform 0 1 2070 -1 0 -4044
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_12
timestamp 1646595912
transform 0 1 2070 -1 0 -4432
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_13
timestamp 1646595912
transform 0 1 2070 -1 0 -4820
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_14
timestamp 1646595912
transform 0 1 2070 -1 0 -5208
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_15
timestamp 1646595912
transform 0 1 2070 -1 0 -5596
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_16
timestamp 1646595912
transform 0 1 2070 -1 0 612
box -224 -2100 224 2100
use sky130_fd_pr__pfet_g5v0d10v5_WL3UED  sky130_fd_pr__pfet_g5v0d10v5_WL3UED_17
timestamp 1646595912
transform 0 1 2070 -1 0 -5984
box -224 -2100 224 2100
use sky130_fd_pr__res_xhigh_po_1p41_P8QAYG  sky130_fd_pr__res_xhigh_po_1p41_P8QAYG_0
timestamp 1725107387
transform 0 1 6342 -1 0 -6093
box -307 -1282 307 1282
<< labels >>
flabel metal1 -1820 3150 -1680 3660 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 -1820 -9510 -1680 -8850 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 8980 1150 9170 2690 0 FreeSans 1600 0 0 0 VOUT
port 3 nsew
flabel metal1 -1820 2370 -1680 2880 0 FreeSans 1600 0 0 0 IB
port 4 nsew
flabel metal1 590 1350 590 1350 0 FreeSans 800 0 0 0 vt
flabel metal2 -350 -6460 -350 -6460 0 FreeSans 800 0 0 0 vl
flabel metal2 4610 -6450 4610 -6450 0 FreeSans 800 0 0 0 vr
flabel metal2 -1820 1130 -1680 1650 0 FreeSans 1600 0 0 0 INN
port 5 nsew
flabel metal2 -1820 -490 -1680 50 0 FreeSans 1600 0 0 0 INP
port 6 nsew
<< properties >>
string MASKHINTS_HVI -1217 -9017 5257 -6583
<< end >>
